module b15s(CK,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G21356,G21357,G21358,G21359,G21360,G21361,G21362,G21363,G21364,G21365,G21366,G21367,G21368,G21369,G21370,G21371,G21372,G21373,G21374,G21375,G21376,G21377,G21378,G21379,G21380,G21381,G21382,G21383,G21384,G21385,G21386,G21387,G21388,G21389,G21794,G21799,G21800,G21802,G21693,G21692,G21691,G21690,G21689,G21688,G21687,G21686,G21685,G21684,G21683,G21682,G21681,G21680,G21679,G21678,G21677,G21676,G21675,G21674,G21673,G21672,G21671,G21670,G21669,G21668,G21667,G21666,G21665,G21664,G21663,G21662);
input CK,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36;
output G21356,G21357,G21358,G21359,G21360,G21361,G21362,G21363,G21364,G21365,G21366,G21367,G21368,G21369,G21370,G21371,G21372,G21373,G21374,G21375,G21376,G21377,G21378,G21379,G21380,G21381,G21382,G21383,G21384,G21385,G21386,G21387,G21388,G21389,G21794,G21799,G21800,G21802,G21693,G21692,G21691,G21690,G21689,G21688,G21687,G21686,G21685,G21684,G21683,G21682,G21681,G21680,G21679,G21678,G21677,G21676,G21675,G21674,G21673,G21672,G21671,G21670,G21669,G21668,G21667,G21666,G21665,G21664,G21663,G21662;

  wire G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
       G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G40,
       G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G60,
       G61,G62,G63,G64,G65,G66,G67,G68,G69,G70,G71,G72,G73,G74,G75,G76,G77,G78,G79,G80,
       G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99,G100,
       G101,G102,G103,G104,G105,G106,G107,G108,G109,G110,G111,G112,G113,G114,G115,G116,G117,G118,G119,G120,
       G121,G122,G123,G124,G125,G126,G127,G128,G129,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G140,
       G141,G142,G143,G144,G145,G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157,G158,G159,G160,
       G161,G162,G163,G164,G165,G166,G167,G168,G169,G170,G171,G172,G173,G174,G175,G176,G177,G178,G179,G180,
       G181,G182,G183,G184,G185,G186,G187,G188,G189,G190,G191,G192,G193,G194,G195,G196,G197,G198,G199,G200,
       G201,G202,G203,G204,G205,G206,G207,G208,G209,G210,G211,G212,G213,G214,G215,G216,G217,G218,G219,G220,
       G221,G222,G223,G224,G225,G226,G227,G228,G229,G230,G231,G232,G233,G234,G235,G236,G237,G238,G239,G240,
       G241,G242,G243,G244,G245,G246,G247,G248,G249,G250,G251,G252,G253,G254,G255,G256,G257,G258,G259,G260,
       G261,G262,G263,G264,G265,G266,G267,G268,G269,G270,G271,G272,G273,G274,G275,G276,G277,G278,G279,G280,
       G281,G282,G283,G284,G285,G286,G287,G288,G289,G290,G291,G292,G293,G294,G295,G296,G297,G298,G299,G300,
       G301,G302,G303,G304,G305,G306,G307,G308,G309,G310,G311,G312,G313,G314,G315,G316,G317,G318,G319,G320,
       G321,G322,G323,G324,G325,G326,G327,G328,G329,G330,G331,G332,G333,G334,G335,G336,G337,G338,G339,G340,
       G341,G342,G343,G344,G345,G346,G347,G348,G349,G350,G351,G352,G353,G354,G355,G356,G357,G358,G359,G360,
       G361,G362,G363,G364,G365,G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,G377,G378,G379,G380,
       G381,G382,G383,G384,G385,G386,G387,G388,G389,G390,G391,G392,G393,G394,G395,G396,G397,G398,G399,G400,
       G401,G402,G403,G404,G405,G406,G407,G408,G409,G410,G411,G412,G413,G414,G415,G416,G417,G418,G419,G420,
       G421,G422,G423,G424,G425,G426,G427,G428,G429,G430,G431,G432,G433,G434,G435,G436,G437,G438,G439,G440,
       G441,G442,G443,G444,G445,G446,G447,G448,G449,G450,G451,G452,G453,G454,G455,G456,G457,G458,G459,G460,
       G461,G462,G463,G464,G465,G466,G467,G468,G469,G470,G471,G472,G473,G474,G475,G476,G477,G478,G479,G480,
       G481,G482,G483,G484,G485,G486,G487,G488,G489,G490,G491,G492,G493,G494,G495,G496,G497,G498,G499,G500,
       G501,G502,G503,G504,G505,G506,G507,G508,G509,G510,G511,G512,G513,G514,G515,G516,G517,G518,G519,G520,
       G521,G522,G523,G524,G525,G526,G527,G528,G529,G530,G531,G532,G533,G534,G535,G536,G537,G538,G539,G540,
       G541,G542,G543,G544,G545,G546,G547,G548,G549,G550,G551,G552,G553,G554,G555,G556,G557,G558,G559,G560,
       G561,G562,G563,G564,G565,G566,G567,G568,G569,G570,G571,G572,G573,G574,G575,G576,G577,G578,G579,G580,
       G581,G582,G583,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G596,G597,G598,G599,G600,
       G601,G602,G603,G604,G605,G606,G607,G608,G609,G610,G611,G612,G613,G614,G615,G616,G617,G618,G619,G620,
       G621,G622,G623,G624,G625,G626,G627,G628,G629,G630,G631,G632,G633,G634,G635,G636,G637,G638,G639,G640,
       G641,G642,G643,G644,G645,G646,G647,G648,G649,G650,G651,G652,G653,G654,G655,G656,G657,G658,G659,G660,
       G661,G662,G663,G664,G665,G666,G667,G668,G669,G670,G671,G672,G673,G674,G675,G676,G677,G678,G679,G680,
       G681,G682,G683,G684,G685,G686,G687,G688,G689,G690,G691,G692,G693,G694,G695,G696,G697,G698,G699,G700,
       G701,G702,G703,G704,G705,G706,G707,G708,G709,G710,G711,G712,G713,G714,G715,G716,G717,G718,G719,G720,
       G721,G722,G723,G724,G725,G726,G727,G728,G729,G730,G731,G732,G733,G734,G735,G736,G737,G738,G739,G740,
       G741,G742,G743,G744,G745,G746,G747,G748,G749,G750,G751,G752,G753,G754,G755,G756,G757,G758,G759,G760,
       G761,G762,G763,G764,G765,G766,G767,G768,G769,G770,G771,G772,G773,G774,G775,G776,G777,G778,G779,G780,
       G781,G782,G783,G784,G785,G786,G787,G788,G789,G790,G791,G792,G793,G794,G795,G796,G797,G798,G799,G800,
       G801,G802,G803,G804,G805,G806,G807,G808,G809,G810,G811,G812,G813,G814,G815,G816,G817,G818,G819,G820,
       G821,G822,G823,G824,G825,G826,G827,G828,G829,G830,G831,G832,G833,G834,G835,G836,G837,G838,G839,G840,
       G841,G842,G843,G844,G845,G846,G847,G848,G849,G850,G851,G852,G853,G854,G855,G856,G857,G858,G859,G860,
       G861,G862,G863,G864,G865,G866,G867,G868,G869,G870,G871,G872,G873,G874,G875,G876,G877,G878,G879,G880,
       G881,G882,G883,G884,G885,G886,G887,G888,G889,G890,G891,G892,G893,G894,G895,G896,G897,G898,G899,G900,
       G901,G902,G903,G904,G905,G906,G907,G908,G909,G910,G911,G912,G913,G914,G915,G916,G917,G918,G919,G920,
       G921,G922,G923,G924,G925,G926,G927,G928,G929,G930,G931,G932,G933,G934,G935,G936,G937,G938,G939,G940,
       G941,G942,G943,G944,G945,G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,G956,G957,G958,G959,G960,
       G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,G971,G972,G973,G974,G975,G976,G977,G978,G979,G980,
       G981,G982,G983,G984,G985,G986,G987,G988,G989,G990,G991,G992,G993,G994,G995,G996,G997,G998,G999,G1000,
       G1001,G1002,G1003,G1004,G1005,G1006,G1007,G1008,G1009,G1010,G1011,G1012,G1013,G1014,G1015,G1016,G1017,G1018,G1019,G1020,
       G1021,G1022,G1023,G1024,G1025,G1026,G1027,G1028,G1029,G1030,G1031,G1032,G1033,G1034,G1035,G1036,G1037,G1038,G1039,G1040,
       G1041,G1042,G1043,G1044,G1045,G1046,G1047,G1048,G1049,G1050,G1051,G1052,G1053,G1054,G1055,G1056,G1057,G1058,G1059,G1060,
       G1061,G1062,G1063,G1064,G1065,G1066,G1067,G1068,G1069,G1070,G1071,G1072,G1073,G1074,G1075,G1076,G1077,G1078,G1079,G1080,
       G1081,G1082,G1083,G1084,G1085,G1086,G1087,G1088,G1089,G1090,G1091,G1092,G1093,G1094,G1095,G1096,G1097,G1098,G1099,G1100,
       G1101,G1102,G1103,G1104,G1105,G1106,G1107,G1108,G1109,G1110,G1111,G1112,G1113,G1114,G1115,G1116,G1117,G1118,G1119,G1120,
       G1121,G1122,G1123,G1124,G1125,G1126,G1127,G1128,G1129,G1130,G1131,G1132,G1133,G1134,G1135,G1136,G1137,G1138,G1139,G1140,
       G1141,G1142,G1143,G1144,G1145,G1146,G1147,G1148,G1149,G1150,G1151,G1152,G1153,G1154,G1155,G1156,G1157,G1158,G1159,G1160,
       G1161,G1162,G1163,G1164,G1165,G1166,G1167,G1168,G1169,G1170,G1171,G1172,G1173,G1174,G1175,G1176,G1177,G1178,G1179,G1180,
       G1181,G1182,G1183,G1184,G1185,G1186,G1187,G1188,G1189,G1190,G1191,G1192,G1193,G1194,G1195,G1196,G1197,G1198,G1199,G1200,
       G1201,G1202,G1203,G1204,G1205,G1206,G1207,G1208,G1209,G1210,G1211,G1212,G1213,G1214,G1215,G1216,G1217,G1218,G1219,G1220,
       G1221,G1222,G1223,G1224,G1225,G1226,G1227,G1228,G1229,G1230,G1231,G1232,G1233,G1234,G1235,G1236,G1237,G1238,G1239,G1240,
       G1241,G1242,G1243,G1244,G1245,G1246,G1247,G1248,G1249,G1250,G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,
       G1261,G1262,G1263,G1264,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272,G1273,G1274,G1275,G1276,G1277,G1278,G1279,G1280,
       G1281,G1282,G1283,G1284,G1285,G1286,G1287,G1288,G1289,G1290,G1291,G1292,G1293,G1294,G1295,G1296,G1297,G1298,G1299,G1300,
       G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,G1310,G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,
       G1321,G1322,G1323,G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,
       G1341,G1342,G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355,G1356,G1357,G1358,G1359,G1360,
       G1361,G1362,G1363,G1364,G1365,G1366,G1367,G1368,G1369,G1370,G1371,G1372,G1373,G1374,G1375,G1376,G1377,G1378,G1379,G1380,
       G1381,G1382,G1383,G1384,G1385,G1386,G1387,G1388,G1389,G1390,G1391,G1392,G1393,G1394,G1395,G1396,G1397,G1398,G1399,G1400,
       G1401,G1402,G1403,G1404,G1405,G1406,G1407,G1408,G1409,G1410,G1411,G1412,G1413,G1414,G1415,G1416,G1417,G1418,G1419,G1420,
       G1421,G1422,G1423,G1424,G1425,G1426,G1427,G1428,G1429,G1430,G1431,G1432,G1433,G1434,G1435,G1436,G1437,G1438,G1439,G1440,
       G1441,G1442,G1443,G1444,G1445,G1446,G1447,G1448,G1449,G1450,G1451,G1452,G1453,G1454,G1455,G1456,G1457,G1458,G1459,G1460,
       G1461,G1462,G1463,G1464,G1465,G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476,G1477,G1478,G1479,G1480,
       G1481,G1482,G1483,G1484,G1485,G1486,G1487,G1488,G1489,G1490,G1491,G1492,G1493,G1494,G1495,G1496,G1497,G1498,G1499,G1500,
       G1501,G1502,G1503,G1504,G1505,G1506,G1507,G1508,G1509,G1510,G1511,G1512,G1513,G1514,G1515,G1516,G1517,G1518,G1519,G1520,
       G1521,G1522,G1523,G1524,G1525,G1526,G1527,G1528,G1529,G1530,G1531,G1532,G1533,G1534,G1535,G1536,G1537,G1538,G1539,G1540,
       G1541,G1542,G1543,G1544,G1545,G1546,G1547,G1548,G1549,G1550,G1551,G1552,G1553,G1554,G1555,G1556,G1557,G1558,G1559,G1560,
       G1561,G1562,G1563,G1564,G1565,G1566,G1567,G1568,G1569,G1570,G1571,G1572,G1573,G1574,G1575,G1576,G1577,G1578,G1579,G1580,
       G1581,G1582,G1583,G1584,G1585,G1586,G1587,G1588,G1589,G1590,G1591,G1592,G1593,G1594,G1595,G1596,G1597,G1598,G1599,G1600,
       G1601,G1602,G1603,G1604,G1605,G1606,G1607,G1608,G1609,G1610,G1611,G1612,G1613,G1614,G1615,G1616,G1617,G1618,G1619,G1620,
       G1621,G1622,G1623,G1624,G1625,G1626,G1627,G1628,G1629,G1630,G1631,G1632,G1633,G1634,G1635,G1636,G1637,G1638,G1639,G1640,
       G1641,G1642,G1643,G1644,G1645,G1646,G1647,G1648,G1649,G1650,G1651,G1652,G1653,G1654,G1655,G1656,G1657,G1658,G1659,G1660,
       G1661,G1662,G1663,G1664,G1665,G1666,G1667,G1668,G1669,G1670,G1671,G1672,G1673,G1674,G1675,G1676,G1677,G1678,G1679,G1680,
       G1681,G1682,G1683,G1684,G1685,G1686,G1687,G1688,G1689,G1690,G1691,G1692,G1693,G1694,G1695,G1696,G1697,G1698,G1699,G1700,
       G1701,G1702,G1703,G1704,G1705,G1706,G1707,G1708,G1709,G1710,G1711,G1712,G1713,G1714,G1715,G1716,G1717,G1718,G1719,G1720,
       G1721,G1722,G1723,G1724,G1725,G1726,G1727,G1728,G1729,G1730,G1731,G1732,G1733,G1734,G1735,G1736,G1737,G1738,G1739,G1740,
       G1741,G1742,G1743,G1744,G1745,G1746,G1747,G1748,G1749,G1750,G1751,G1752,G1753,G1754,G1755,G1756,G1757,G1758,G1759,G1760,
       G1761,G1762,G1763,G1764,G1765,G1766,G1767,G1768,G1769,G1770,G1771,G1772,G1773,G1774,G1775,G1776,G1777,G1778,G1779,G1780,
       G1781,G1782,G1783,G1784,G1785,G1786,G1787,G1788,G1789,G1790,G1791,G1792,G1793,G1794,G1795,G1796,G1797,G1798,G1799,G1800,
       G1801,G1802,G1803,G1804,G1805,G1806,G1807,G1808,G1809,G1810,G1811,G1812,G1813,G1814,G1815,G1816,G1817,G1818,G1819,G1820,
       G1821,G1822,G1823,G1824,G1825,G1826,G1827,G1828,G1829,G1830,G1831,G1832,G1833,G1834,G1835,G1836,G1837,G1838,G1839,G1840,
       G1841,G1842,G1843,G1844,G1845,G1846,G1847,G1848,G1849,G1850,G1851,G1852,G1853,G1854,G1855,G1856,G1857,G1858,G1859,G1860,
       G1861,G1862,G1863,G1864,G1865,G1866,G1867,G1868,G1869,G1870,G1871,G1872,G1873,G1874,G1875,G1876,G1877,G1878,G1879,G1880,
       G1881,G1882,G1883,G1884,G1885,G1886,G1887,G1888,G1889,G1890,G1891,G1892,G1893,G1894,G1895,G1896,G1897,G1898,G1899,G1900,
       G1901,G1902,G1903,G1904,G1905,G1906,G1907,G1908,G1909,G1910,G1911,G1912,G1913,G1914,G1915,G1916,G1917,G1918,G1919,G1920,
       G1921,G1922,G1923,G1924,G1925,G1926,G1927,G1928,G1929,G1930,G1931,G1932,G1933,G1934,G1935,G1936,G1937,G1938,G1939,G1940,
       G1941,G1942,G1943,G1944,G1945,G1946,G1947,G1948,G1949,G1950,G1951,G1952,G1953,G1954,G1955,G1956,G1957,G1958,G1959,G1960,
       G1961,G1962,G1963,G1964,G1965,G1966,G1967,G1968,G1969,G1970,G1971,G1972,G1973,G1974,G1975,G1976,G1977,G1978,G1979,G1980,
       G1981,G1982,G1983,G1984,G1985,G1986,G1987,G1988,G1989,G1990,G1991,G1992,G1993,G1994,G1995,G1996,G1997,G1998,G1999,G2000,
       G2001,G2002,G2003,G2004,G2005,G2006,G2007,G2008,G2009,G2010,G2011,G2012,G2013,G2014,G2015,G2016,G2017,G2018,G2019,G2020,
       G2021,G2022,G2023,G2024,G2025,G2026,G2027,G2028,G2029,G2030,G2031,G2032,G2033,G2034,G2035,G2036,G2037,G2038,G2039,G2040,
       G2041,G2042,G2043,G2044,G2045,G2046,G2047,G2048,G2049,G2050,G2051,G2052,G2053,G2054,G2055,G2056,G2057,G2058,G2059,G2060,
       G2061,G2062,G2063,G2064,G2065,G2066,G2067,G2068,G2069,G2070,G2071,G2072,G2073,G2074,G2075,G2076,G2077,G2078,G2079,G2080,
       G2081,G2082,G2083,G2084,G2085,G2086,G2087,G2088,G2089,G2090,G2091,G2092,G2093,G2094,G2095,G2096,G2097,G2098,G2099,G2100,
       G2101,G2102,G2103,G2104,G2105,G2106,G2107,G2108,G2109,G2110,G2111,G2112,G2113,G2114,G2115,G2116,G2117,G2118,G2119,G2120,
       G2121,G2122,G2123,G2124,G2125,G2126,G2127,G2128,G2129,G2130,G2131,G2132,G2133,G2134,G2135,G2136,G2137,G2138,G2139,G2140,
       G2141,G2142,G2143,G2144,G2145,G2146,G2147,G2148,G2149,G2150,G2151,G2152,G2153,G2154,G2155,G2156,G2157,G2158,G2159,G2160,
       G2161,G2162,G2163,G2164,G2165,G2166,G2167,G2168,G2169,G2170,G2171,G2172,G2173,G2174,G2175,G2176,G2177,G2178,G2179,G2180,
       G2181,G2182,G2183,G2184,G2185,G2186,G2187,G2188,G2189,G2190,G2191,G2192,G2193,G2194,G2195,G2196,G2197,G2198,G2199,G2200,
       G2201,G2202,G2203,G2204,G2205,G2206,G2207,G2208,G2209,G2210,G2211,G2212,G2213,G2214,G2215,G2216,G2217,G2218,G2219,G2220,
       G2221,G2222,G2223,G2224,G2225,G2226,G2227,G2228,G2229,G2230,G2231,G2232,G2233,G2234,G2235,G2236,G2237,G2238,G2239,G2240,
       G2241,G2242,G2243,G2244,G2245,G2246,G2247,G2248,G2249,G2250,G2251,G2252,G2253,G2254,G2255,G2256,G2257,G2258,G2259,G2260,
       G2261,G2262,G2263,G2264,G2265,G2266,G2267,G2268,G2269,G2270,G2271,G2272,G2273,G2274,G2275,G2276,G2277,G2278,G2279,G2280,
       G2281,G2282,G2283,G2284,G2285,G2286,G2287,G2288,G2289,G2290,G2291,G2292,G2293,G2294,G2295,G2296,G2297,G2298,G2299,G2300,
       G2301,G2302,G2303,G2304,G2305,G2306,G2307,G2308,G2309,G2310,G2311,G2312,G2313,G2314,G2315,G2316,G2317,G2318,G2319,G2320,
       G2321,G2322,G2323,G2324,G2325,G2326,G2327,G2328,G2329,G2330,G2331,G2332,G2333,G2334,G2335,G2336,G2337,G2338,G2339,G2340,
       G2341,G2342,G2343,G2344,G2345,G2346,G2347,G2348,G2349,G2350,G2351,G2352,G2353,G2354,G2355,G2356,G2357,G2358,G2359,G2360,
       G2361,G2362,G2363,G2364,G2365,G2366,G2367,G2368,G2369,G2370,G2371,G2372,G2373,G2374,G2375,G2376,G2377,G2378,G2379,G2380,
       G2381,G2382,G2383,G2384,G2385,G2386,G2387,G2388,G2389,G2390,G2391,G2392,G2393,G2394,G2395,G2396,G2397,G2398,G2399,G2400,
       G2401,G2402,G2403,G2404,G2405,G2406,G2407,G2408,G2409,G2410,G2411,G2412,G2413,G2414,G2415,G2416,G2417,G2418,G2419,G2420,
       G2421,G2422,G2423,G2424,G2425,G2426,G2427,G2428,G2429,G2430,G2431,G2432,G2433,G2434,G2435,G2436,G2437,G2438,G2439,G2440,
       G2441,G2442,G2443,G2444,G2445,G2446,G2447,G2448,G2449,G2450,G2451,G2452,G2453,G2454,G2455,G2456,G2457,G2458,G2459,G2460,
       G2461,G2462,G2463,G2464,G2465,G2466,G2467,G2468,G2469,G2470,G2471,G2472,G2473,G2474,G2475,G2476,G2477,G2478,G2479,G2480,
       G2481,G2482,G2483,G2484,G2485,G2486,G2487,G2488,G2489,G2490,G2491,G2492,G2493,G2494,G2495,G2496,G2497,G2498,G2499,G2500,
       G2501,G2502,G2503,G2504,G2505,G2506,G2507,G2508,G2509,G2510,G2511,G2512,G2513,G2514,G2515,G2516,G2517,G2518,G2519,G2520,
       G2521,G2522,G2523,G2524,G2525,G2526,G2527,G2528,G2529,G2530,G2531,G2532,G2533,G2534,G2535,G2536,G2537,G2538,G2539,G2540,
       G2541,G2542,G2543,G2544,G2545,G2546,G2547,G2548,G2549,G2550,G2551,G2552,G2553,G2554,G2555,G2556,G2557,G2558,G2559,G2560,
       G2561,G2562,G2563,G2564,G2565,G2566,G2567,G2568,G2569,G2570,G2571,G2572,G2573,G2574,G2575,G2576,G2577,G2578,G2579,G2580,
       G2581,G2582,G2583,G2584,G2585,G2586,G2587,G2588,G2589,G2590,G2591,G2592,G2593,G2594,G2595,G2596,G2597,G2598,G2599,G2600,
       G2601,G2602,G2603,G2604,G2605,G2606,G2607,G2608,G2609,G2610,G2611,G2612,G2613,G2614,G2615,G2616,G2617,G2618,G2619,G2620,
       G2621,G2622,G2623,G2624,G2625,G2626,G2627,G2628,G2629,G2630,G2631,G2632,G2633,G2634,G2635,G2636,G2637,G2638,G2639,G2640,
       G2641,G2642,G2643,G2644,G2645,G2646,G2647,G2648,G2649,G2650,G2651,G2652,G2653,G2654,G2655,G2656,G2657,G2658,G2659,G2660,
       G2661,G2662,G2663,G2664,G2665,G2666,G2667,G2668,G2669,G2670,G2671,G2672,G2673,G2674,G2675,G2676,G2677,G2678,G2679,G2680,
       G2681,G2682,G2683,G2684,G2685,G2686,G2687,G2688,G2689,G2690,G2691,G2692,G2693,G2694,G2695,G2696,G2697,G2698,G2699,G2700,
       G2701,G2702,G2703,G2704,G2705,G2706,G2707,G2708,G2709,G2710,G2711,G2712,G2713,G2714,G2715,G2716,G2717,G2718,G2719,G2720,
       G2721,G2722,G2723,G2724,G2725,G2726,G2727,G2728,G2729,G2730,G2731,G2732,G2733,G2734,G2735,G2736,G2737,G2738,G2739,G2740,
       G2741,G2742,G2743,G2744,G2745,G2746,G2747,G2748,G2749,G2750,G2751,G2752,G2753,G2754,G2755,G2756,G2757,G2758,G2759,G2760,
       G2761,G2762,G2763,G2764,G2765,G2766,G2767,G2768,G2769,G2770,G2771,G2772,G2773,G2774,G2775,G2776,G2777,G2778,G2779,G2780,
       G2781,G2782,G2783,G2784,G2785,G2786,G2787,G2788,G2789,G2790,G2791,G2792,G2793,G2794,G2795,G2796,G2797,G2798,G2799,G2800,
       G2801,G2802,G2803,G2804,G2805,G2806,G2807,G2808,G2809,G2810,G2811,G2812,G2813,G2814,G2815,G2816,G2817,G2818,G2819,G2820,
       G2821,G2822,G2823,G2824,G2825,G2826,G2827,G2828,G2829,G2830,G2831,G2832,G2833,G2834,G2835,G2836,G2837,G2838,G2839,G2840,
       G2841,G2842,G2843,G2844,G2845,G2846,G2847,G2848,G2849,G2850,G2851,G2852,G2853,G2854,G2855,G2856,G2857,G2858,G2859,G2860,
       G2861,G2862,G2863,G2864,G2865,G2866,G2867,G2868,G2869,G2870,G2871,G2872,G2873,G2874,G2875,G2876,G2877,G2878,G2879,G2880,
       G2881,G2882,G2883,G2884,G2885,G2886,G2887,G2888,G2889,G2890,G2891,G2892,G2893,G2894,G2895,G2896,G2897,G2898,G2899,G2900,
       G2901,G2902,G2903,G2904,G2905,G2906,G2907,G2908,G2909,G2910,G2911,G2912,G2913,G2914,G2915,G2916,G2917,G2918,G2919,G2920,
       G2921,G2922,G2923,G2924,G2925,G2926,G2927,G2928,G2929,G2930,G2931,G2932,G2933,G2934,G2935,G2936,G2937,G2938,G2939,G2940,
       G2941,G2942,G2943,G2944,G2945,G2946,G2947,G2948,G2949,G2950,G2951,G2952,G2953,G2954,G2955,G2956,G2957,G2958,G2959,G2960,
       G2961,G2962,G2963,G2964,G2965,G2966,G2967,G2968,G2969,G2970,G2971,G2972,G2973,G2974,G2975,G2976,G2977,G2978,G2979,G2980,
       G2981,G2982,G2983,G2984,G2985,G2986,G2987,G2988,G2989,G2990,G2991,G2992,G2993,G2994,G2995,G2996,G2997,G2998,G2999,G3000,
       G3001,G3002,G3003,G3004,G3005,G3006,G3007,G3008,G3009,G3010,G3011,G3012,G3013,G3014,G3015,G3016,G3017,G3018,G3019,G3020,
       G3021,G3022,G3023,G3024,G3025,G3026,G3027,G3028,G3029,G3030,G3031,G3032,G3033,G3034,G3035,G3036,G3037,G3038,G3039,G3040,
       G3041,G3042,G3043,G3044,G3045,G3046,G3047,G3048,G3049,G3050,G3051,G3052,G3053,G3054,G3055,G3056,G3057,G3058,G3059,G3060,
       G3061,G3062,G3063,G3064,G3065,G3066,G3067,G3068,G3069,G3070,G3071,G3072,G3073,G3074,G3075,G3076,G3077,G3078,G3079,G3080,
       G3081,G3082,G3083,G3084,G3085,G3086,G3087,G3088,G3089,G3090,G3091,G3092,G3093,G3094,G3095,G3096,G3097,G3098,G3099,G3100,
       G3101,G3102,G3103,G3104,G3105,G3106,G3107,G3108,G3109,G3110,G3111,G3112,G3113,G3114,G3115,G3116,G3117,G3118,G3119,G3120,
       G3121,G3122,G3123,G3124,G3125,G3126,G3127,G3128,G3129,G3130,G3131,G3132,G3133,G3134,G3135,G3136,G3137,G3138,G3139,G3140,
       G3141,G3142,G3143,G3144,G3145,G3146,G3147,G3148,G3149,G3150,G3151,G3152,G3153,G3154,G3155,G3156,G3157,G3158,G3159,G3160,
       G3161,G3162,G3163,G3164,G3165,G3166,G3167,G3168,G3169,G3170,G3171,G3172,G3173,G3174,G3175,G3176,G3177,G3178,G3179,G3180,
       G3181,G3182,G3183,G3184,G3185,G3186,G3187,G3188,G3189,G3190,G3191,G3192,G3193,G3194,G3195,G3196,G3197,G3198,G3199,G3200,
       G3201,G3202,G3203,G3204,G3205,G3206,G3207,G3208,G3209,G3210,G3211,G3212,G3213,G3214,G3215,G3216,G3217,G3218,G3219,G3220,
       G3221,G3222,G3223,G3224,G3225,G3226,G3227,G3228,G3229,G3230,G3231,G3232,G3233,G3234,G3235,G3236,G3237,G3238,G3239,G3240,
       G3241,G3242,G3243,G3244,G3245,G3246,G3247,G3248,G3249,G3250,G3251,G3252,G3253,G3254,G3255,G3256,G3257,G3258,G3259,G3260,
       G3261,G3262,G3263,G3264,G3265,G3266,G3267,G3268,G3269,G3270,G3271,G3272,G3273,G3274,G3275,G3276,G3277,G3278,G3279,G3280,
       G3281,G3282,G3283,G3284,G3285,G3286,G3287,G3288,G3289,G3290,G3291,G3292,G3293,G3294,G3295,G3296,G3297,G3298,G3299,G3300,
       G3301,G3302,G3303,G3304,G3305,G3306,G3307,G3308,G3309,G3310,G3311,G3312,G3313,G3314,G3315,G3316,G3317,G3318,G3319,G3320,
       G3321,G3322,G3323,G3324,G3325,G3326,G3327,G3328,G3329,G3330,G3331,G3332,G3333,G3334,G3335,G3336,G3337,G3338,G3339,G3340,
       G3341,G3342,G3343,G3344,G3345,G3346,G3347,G3348,G3349,G3350,G3351,G3352,G3353,G3354,G3355,G3356,G3357,G3358,G3359,G3360,
       G3361,G3362,G3363,G3364,G3365,G3366,G3367,G3368,G3369,G3370,G3371,G3372,G3373,G3374,G3375,G3376,G3377,G3378,G3379,G3380,
       G3381,G3382,G3383,G3384,G3385,G3386,G3387,G3388,G3389,G3390,G3391,G3392,G3393,G3394,G3395,G3396,G3397,G3398,G3399,G3400,
       G3401,G3402,G3403,G3404,G3405,G3406,G3407,G3408,G3409,G3410,G3411,G3412,G3413,G3414,G3415,G3416,G3417,G3418,G3419,G3420,
       G3421,G3422,G3423,G3424,G3425,G3426,G3427,G3428,G3429,G3430,G3431,G3432,G3433,G3434,G3435,G3436,G3437,G3438,G3439,G3440,
       G3441,G3442,G3443,G3444,G3445,G3446,G3447,G3448,G3449,G3450,G3451,G3452,G3453,G3454,G3455,G3456,G3457,G3458,G3459,G3460,
       G3461,G3462,G3463,G3464,G3465,G3466,G3467,G3468,G3469,G3470,G3471,G3472,G3473,G3474,G3475,G3476,G3477,G3478,G3479,G3480,
       G3481,G3482,G3483,G3484,G3485,G3486,G3487,G3488,G3489,G3490,G3491,G3492,G3493,G3494,G3495,G3496,G3497,G3498,G3499,G3500,
       G3501,G3502,G3503,G3504,G3505,G3506,G3507,G3508,G3509,G3510,G3511,G3512,G3513,G3514,G3515,G3516,G3517,G3518,G3519,G3520,
       G3521,G3522,G3523,G3524,G3525,G3526,G3527,G3528,G3529,G3530,G3531,G3532,G3533,G3534,G3535,G3536,G3537,G3538,G3539,G3540,
       G3541,G3542,G3543,G3544,G3545,G3546,G3547,G3548,G3549,G3550,G3551,G3552,G3553,G3554,G3555,G3556,G3557,G3558,G3559,G3560,
       G3561,G3562,G3563,G3564,G3565,G3566,G3567,G3568,G3569,G3570,G3571,G3572,G3573,G3574,G3575,G3576,G3577,G3578,G3579,G3580,
       G3581,G3582,G3583,G3584,G3585,G3586,G3587,G3588,G3589,G3590,G3591,G3592,G3593,G3594,G3595,G3596,G3597,G3598,G3599,G3600,
       G3601,G3602,G3603,G3604,G3605,G3606,G3607,G3608,G3609,G3610,G3611,G3612,G3613,G3614,G3615,G3616,G3617,G3618,G3619,G3620,
       G3621,G3622,G3623,G3624,G3625,G3626,G3627,G3628,G3629,G3630,G3631,G3632,G3633,G3634,G3635,G3636,G3637,G3638,G3639,G3640,
       G3641,G3642,G3643,G3644,G3645,G3646,G3647,G3648,G3649,G3650,G3651,G3652,G3653,G3654,G3655,G3656,G3657,G3658,G3659,G3660,
       G3661,G3662,G3663,G3664,G3665,G3666,G3667,G3668,G3669,G3670,G3671,G3672,G3673,G3674,G3675,G3676,G3677,G3678,G3679,G3680,
       G3681,G3682,G3683,G3684,G3685,G3686,G3687,G3688,G3689,G3690,G3691,G3692,G3693,G3694,G3695,G3696,G3697,G3698,G3699,G3700,
       G3701,G3702,G3703,G3704,G3705,G3706,G3707,G3708,G3709,G3710,G3711,G3712,G3713,G3714,G3715,G3716,G3717,G3718,G3719,G3720,
       G3721,G3722,G3723,G3724,G3725,G3726,G3727,G3728,G3729,G3730,G3731,G3732,G3733,G3734,G3735,G3736,G3737,G3738,G3739,G3740,
       G3741,G3742,G3743,G3744,G3745,G3746,G3747,G3748,G3749,G3750,G3751,G3752,G3753,G3754,G3755,G3756,G3757,G3758,G3759,G3760,
       G3761,G3762,G3763,G3764,G3765,G3766,G3767,G3768,G3769,G3770,G3771,G3772,G3773,G3774,G3775,G3776,G3777,G3778,G3779,G3780,
       G3781,G3782,G3783,G3784,G3785,G3786,G3787,G3788,G3789,G3790,G3791,G3792,G3793,G3794,G3795,G3796,G3797,G3798,G3799,G3800,
       G3801,G3802,G3803,G3804,G3805,G3806,G3807,G3808,G3809,G3810,G3811,G3812,G3813,G3814,G3815,G3816,G3817,G3818,G3819,G3820,
       G3821,G3822,G3823,G3824,G3825,G3826,G3827,G3828,G3829,G3830,G3831,G3832,G3833,G3834,G3835,G3836,G3837,G3838,G3839,G3840,
       G3841,G3842,G3843,G3844,G3845,G3846,G3847,G3848,G3849,G3850,G3851,G3852,G3853,G3854,G3855,G3856,G3857,G3858,G3859,G3860,
       G3861,G3862,G3863,G3864,G3865,G3866,G3867,G3868,G3869,G3870,G3871,G3872,G3873,G3874,G3875,G3876,G3877,G3878,G3879,G3880,
       G3881,G3882,G3883,G3884,G3885,G3886,G3887,G3888,G3889,G3890,G3891,G3892,G3893,G3894,G3895,G3896,G3897,G3898,G3899,G3900,
       G3901,G3902,G3903,G3904,G3905,G3906,G3907,G3908,G3909,G3910,G3911,G3912,G3913,G3914,G3915,G3916,G3917,G3918,G3919,G3920,
       G3921,G3922,G3923,G3924,G3925,G3926,G3927,G3928,G3929,G3930,G3931,G3932,G3933,G3934,G3935,G3936,G3937,G3938,G3939,G3940,
       G3941,G3942,G3943,G3944,G3945,G3946,G3947,G3948,G3949,G3950,G3951,G3952,G3953,G3954,G3955,G3956,G3957,G3958,G3959,G3960,
       G3961,G3962,G3963,G3964,G3965,G3966,G3967,G3968,G3969,G3970,G3971,G3972,G3973,G3974,G3975,G3976,G3977,G3978,G3979,G3980,
       G3981,G3982,G3983,G3984,G3985,G3986,G3987,G3988,G3989,G3990,G3991,G3992,G3993,G3994,G3995,G3996,G3997,G3998,G3999,G4000,
       G4001,G4002,G4003,G4004,G4005,G4006,G4007,G4008,G4009,G4010,G4011,G4012,G4013,G4014,G4015,G4016,G4017,G4018,G4019,G4020,
       G4021,G4022,G4023,G4024,G4025,G4026,G4027,G4028,G4029,G4030,G4031,G4032,G4033,G4034,G4035,G4036,G4037,G4038,G4039,G4040,
       G4041,G4042,G4043,G4044,G4045,G4046,G4047,G4048,G4049,G4050,G4051,G4052,G4053,G4054,G4055,G4056,G4057,G4058,G4059,G4060,
       G4061,G4062,G4063,G4064,G4065,G4066,G4067,G4068,G4069,G4070,G4071,G4072,G4073,G4074,G4075,G4076,G4077,G4078,G4079,G4080,
       G4081,G4082,G4083,G4084,G4085,G4086,G4087,G4088,G4089,G4090,G4091,G4092,G4093,G4094,G4095,G4096,G4097,G4098,G4099,G4100,
       G4101,G4102,G4103,G4104,G4105,G4106,G4107,G4108,G4109,G4110,G4111,G4112,G4113,G4114,G4115,G4116,G4117,G4118,G4119,G4120,
       G4121,G4122,G4123,G4124,G4125,G4126,G4127,G4128,G4129,G4130,G4131,G4132,G4133,G4134,G4135,G4136,G4137,G4138,G4139,G4140,
       G4141,G4142,G4143,G4144,G4145,G4146,G4147,G4148,G4149,G4150,G4151,G4152,G4153,G4154,G4155,G4156,G4157,G4158,G4159,G4160,
       G4161,G4162,G4163,G4164,G4165,G4166,G4167,G4168,G4169,G4170,G4171,G4172,G4173,G4174,G4175,G4176,G4177,G4178,G4179,G4180,
       G4181,G4182,G4183,G4184,G4185,G4186,G4187,G4188,G4189,G4190,G4191,G4192,G4193,G4194,G4195,G4196,G4197,G4198,G4199,G4200,
       G4201,G4202,G4203,G4204,G4205,G4206,G4207,G4208,G4209,G4210,G4211,G4212,G4213,G4214,G4215,G4216,G4217,G4218,G4219,G4220,
       G4221,G4222,G4223,G4224,G4225,G4226,G4227,G4228,G4229,G4230,G4231,G4232,G4233,G4234,G4235,G4236,G4237,G4238,G4239,G4240,
       G4241,G4242,G4243,G4244,G4245,G4246,G4247,G4248,G4249,G4250,G4251,G4252,G4253,G4254,G4255,G4256,G4257,G4258,G4259,G4260,
       G4261,G4262,G4263,G4264,G4265,G4266,G4267,G4268,G4269,G4270,G4271,G4272,G4273,G4274,G4275,G4276,G4277,G4278,G4279,G4280,
       G4281,G4282,G4283,G4284,G4285,G4286,G4287,G4288,G4289,G4290,G4291,G4292,G4293,G4294,G4295,G4296,G4297,G4298,G4299,G4300,
       G4301,G4302,G4303,G4304,G4305,G4306,G4307,G4308,G4309,G4310,G4311,G4312,G4313,G4314,G4315,G4316,G4317,G4318,G4319,G4320,
       G4321,G4322,G4323,G4324,G4325,G4326,G4327,G4328,G4329,G4330,G4331,G4332,G4333,G4334,G4335,G4336,G4337,G4338,G4339,G4340,
       G4341,G4342,G4343,G4344,G4345,G4346,G4347,G4348,G4349,G4350,G4351,G4352,G4353,G4354,G4355,G4356,G4357,G4358,G4359,G4360,
       G4361,G4362,G4363,G4364,G4365,G4366,G4367,G4368,G4369,G4370,G4371,G4372,G4373,G4374,G4375,G4376,G4377,G4378,G4379,G4380,
       G4381,G4382,G4383,G4384,G4385,G4386,G4387,G4388,G4389,G4390,G4391,G4392,G4393,G4394,G4395,G4396,G4397,G4398,G4399,G4400,
       G4401,G4402,G4403,G4404,G4405,G4406,G4407,G4408,G4409,G4410,G4411,G4412,G4413,G4414,G4415,G4416,G4417,G4418,G4419,G4420,
       G4421,G4422,G4423,G4424,G4425,G4426,G4427,G4428,G4429,G4430,G4431,G4432,G4433,G4434,G4435,G4436,G4437,G4438,G4439,G4440,
       G4441,G4442,G4443,G4444,G4445,G4446,G4447,G4448,G4449,G4450,G4451,G4452,G4453,G4454,G4455,G4456,G4457,G4458,G4459,G4460,
       G4461,G4462,G4463,G4464,G4465,G4466,G4467,G4468,G4469,G4470,G4471,G4472,G4473,G4474,G4475,G4476,G4477,G4478,G4479,G4480,
       G4481,G4482,G4483,G4484,G4485,G4486,G4487,G4488,G4489,G4490,G4491,G4492,G4493,G4494,G4495,G4496,G4497,G4498,G4499,G4500,
       G4501,G4502,G4503,G4504,G4505,G4506,G4507,G4508,G4509,G4510,G4511,G4512,G4513,G4514,G4515,G4516,G4517,G4518,G4519,G4520,
       G4521,G4522,G4523,G4524,G4525,G4526,G4527,G4528,G4529,G4530,G4531,G4532,G4533,G4534,G4535,G4536,G4537,G4538,G4539,G4540,
       G4541,G4542,G4543,G4544,G4545,G4546,G4547,G4548,G4549,G4550,G4551,G4552,G4553,G4554,G4555,G4556,G4557,G4558,G4559,G4560,
       G4561,G4562,G4563,G4564,G4565,G4566,G4567,G4568,G4569,G4570,G4571,G4572,G4573,G4574,G4575,G4576,G4577,G4578,G4579,G4580,
       G4581,G4582,G4583,G4584,G4585,G4586,G4587,G4588,G4589,G4590,G4591,G4592,G4593,G4594,G4595,G4596,G4597,G4598,G4599,G4600,
       G4601,G4602,G4603,G4604,G4605,G4606,G4607,G4608,G4609,G4610,G4611,G4612,G4613,G4614,G4615,G4616,G4617,G4618,G4619,G4620,
       G4621,G4622,G4623,G4624,G4625,G4626,G4627,G4628,G4629,G4630,G4631,G4632,G4633,G4634,G4635,G4636,G4637,G4638,G4639,G4640,
       G4641,G4642,G4643,G4644,G4645,G4646,G4647,G4648,G4649,G4650,G4651,G4652,G4653,G4654,G4655,G4656,G4657,G4658,G4659,G4660,
       G4661,G4662,G4663,G4664,G4665,G4666,G4667,G4668,G4669,G4670,G4671,G4672,G4673,G4674,G4675,G4676,G4677,G4678,G4679,G4680,
       G4681,G4682,G4683,G4684,G4685,G4686,G4687,G4688,G4689,G4690,G4691,G4692,G4693,G4694,G4695,G4696,G4697,G4698,G4699,G4700,
       G4701,G4702,G4703,G4704,G4705,G4706,G4707,G4708,G4709,G4710,G4711,G4712,G4713,G4714,G4715,G4716,G4717,G4718,G4719,G4720,
       G4721,G4722,G4723,G4724,G4725,G4726,G4727,G4728,G4729,G4730,G4731,G4732,G4733,G4734,G4735,G4736,G4737,G4738,G4739,G4740,
       G4741,G4742,G4743,G4744,G4745,G4746,G4747,G4748,G4749,G4750,G4751,G4752,G4753,G4754,G4755,G4756,G4757,G4758,G4759,G4760,
       G4761,G4762,G4763,G4764,G4765,G4766,G4767,G4768,G4769,G4770,G4771,G4772,G4773,G4774,G4775,G4776,G4777,G4778,G4779,G4780,
       G4781,G4782,G4783,G4784,G4785,G4786,G4787,G4788,G4789,G4790,G4791,G4792,G4793,G4794,G4795,G4796,G4797,G4798,G4799,G4800,
       G4801,G4802,G4803,G4804,G4805,G4806,G4807,G4808,G4809,G4810,G4811,G4812,G4813,G4814,G4815,G4816,G4817,G4818,G4819,G4820,
       G4821,G4822,G4823,G4824,G4825,G4826,G4827,G4828,G4829,G4830,G4831,G4832,G4833,G4834,G4835,G4836,G4837,G4838,G4839,G4840,
       G4841,G4842,G4843,G4844,G4845,G4846,G4847,G4848,G4849,G4850,G4851,G4852,G4853,G4854,G4855,G4856,G4857,G4858,G4859,G4860,
       G4861,G4862,G4863,G4864,G4865,G4866,G4867,G4868,G4869,G4870,G4871,G4872,G4873,G4874,G4875,G4876,G4877,G4878,G4879,G4880,
       G4881,G4882,G4883,G4884,G4885,G4886,G4887,G4888,G4889,G4890,G4891,G4892,G4893,G4894,G4895,G4896,G4897,G4898,G4899,G4900,
       G4901,G4902,G4903,G4904,G4905,G4906,G4907,G4908,G4909,G4910,G4911,G4912,G4913,G4914,G4915,G4916,G4917,G4918,G4919,G4920,
       G4921,G4922,G4923,G4924,G4925,G4926,G4927,G4928,G4929,G4930,G4931,G4932,G4933,G4934,G4935,G4936,G4937,G4938,G4939,G4940,
       G4941,G4942,G4943,G4944,G4945,G4946,G4947,G4948,G4949,G4950,G4951,G4952,G4953,G4954,G4955,G4956,G4957,G4958,G4959,G4960,
       G4961,G4962,G4963,G4964,G4965,G4966,G4967,G4968,G4969,G4970,G4971,G4972,G4973,G4974,G4975,G4976,G4977,G4978,G4979,G4980,
       G4981,G4982,G4983,G4984,G4985,G4986,G4987,G4988,G4989,G4990,G4991,G4992,G4993,G4994,G4995,G4996,G4997,G4998,G4999,G5000,
       G5001,G5002,G5003,G5004,G5005,G5006,G5007,G5008,G5009,G5010,G5011,G5012,G5013,G5014,G5015,G5016,G5017,G5018,G5019,G5020,
       G5021,G5022,G5023,G5024,G5025,G5026,G5027,G5028,G5029,G5030,G5031,G5032,G5033,G5034,G5035,G5036,G5037,G5038,G5039,G5040,
       G5041,G5042,G5043,G5044,G5045,G5046,G5047,G5048,G5049,G5050,G5051,G5052,G5053,G5054,G5055,G5056,G5057,G5058,G5059,G5060,
       G5061,G5062,G5063,G5064,G5065,G5066,G5067,G5068,G5069,G5070,G5071,G5072,G5073,G5074,G5075,G5076,G5077,G5078,G5079,G5080,
       G5081,G5082,G5083,G5084,G5085,G5086,G5087,G5088,G5089,G5090,G5091,G5092,G5093,G5094,G5095,G5096,G5097,G5098,G5099,G5100,
       G5101,G5102,G5103,G5104,G5105,G5106,G5107,G5108,G5109,G5110,G5111,G5112,G5113,G5114,G5115,G5116,G5117,G5118,G5119,G5120,
       G5121,G5122,G5123,G5124,G5125,G5126,G5127,G5128,G5129,G5130,G5131,G5132,G5133,G5134,G5135,G5136,G5137,G5138,G5139,G5140,
       G5141,G5142,G5143,G5144,G5145,G5146,G5147,G5148,G5149,G5150,G5151,G5152,G5153,G5154,G5155,G5156,G5157,G5158,G5159,G5160,
       G5161,G5162,G5163,G5164,G5165,G5166,G5167,G5168,G5169,G5170,G5171,G5172,G5173,G5174,G5175,G5176,G5177,G5178,G5179,G5180,
       G5181,G5182,G5183,G5184,G5185,G5186,G5187,G5188,G5189,G5190,G5191,G5192,G5193,G5194,G5195,G5196,G5197,G5198,G5199,G5200,
       G5201,G5202,G5203,G5204,G5205,G5206,G5207,G5208,G5209,G5210,G5211,G5212,G5213,G5214,G5215,G5216,G5217,G5218,G5219,G5220,
       G5221,G5222,G5223,G5224,G5225,G5226,G5227,G5228,G5229,G5230,G5231,G5232,G5233,G5234,G5235,G5236,G5237,G5238,G5239,G5240,
       G5241,G5242,G5243,G5244,G5245,G5246,G5247,G5248,G5249,G5250,G5251,G5252,G5253,G5254,G5255,G5256,G5257,G5258,G5259,G5260,
       G5261,G5262,G5263,G5264,G5265,G5266,G5267,G5268,G5269,G5270,G5271,G5272,G5273,G5274,G5275,G5276,G5277,G5278,G5279,G5280,
       G5281,G5282,G5283,G5284,G5285,G5286,G5287,G5288,G5289,G5290,G5291,G5292,G5293,G5294,G5295,G5296,G5297,G5298,G5299,G5300,
       G5301,G5302,G5303,G5304,G5305,G5306,G5307,G5308,G5309,G5310,G5311,G5312,G5313,G5314,G5315,G5316,G5317,G5318,G5319,G5320,
       G5321,G5322,G5323,G5324,G5325,G5326,G5327,G5328,G5329,G5330,G5331,G5332,G5333,G5334,G5335,G5336,G5337,G5338,G5339,G5340,
       G5341,G5342,G5343,G5344,G5345,G5346,G5347,G5348,G5349,G5350,G5351,G5352,G5353,G5354,G5355,G5356,G5357,G5358,G5359,G5360,
       G5361,G5362,G5363,G5364,G5365,G5366,G5367,G5368,G5369,G5370,G5371,G5372,G5373,G5374,G5375,G5376,G5377,G5378,G5379,G5380,
       G5381,G5382,G5383,G5384,G5385,G5386,G5387,G5388,G5389,G5390,G5391,G5392,G5393,G5394,G5395,G5396,G5397,G5398,G5399,G5400,
       G5401,G5402,G5403,G5404,G5405,G5406,G5407,G5408,G5409,G5410,G5411,G5412,G5413,G5414,G5415,G5416,G5417,G5418,G5419,G5420,
       G5421,G5422,G5423,G5424,G5425,G5426,G5427,G5428,G5429,G5430,G5431,G5432,G5433,G5434,G5435,G5436,G5437,G5438,G5439,G5440,
       G5441,G5442,G5443,G5444,G5445,G5446,G5447,G5448,G5449,G5450,G5451,G5452,G5453,G5454,G5455,G5456,G5457,G5458,G5459,G5460,
       G5461,G5462,G5463,G5464,G5465,G5466,G5467,G5468,G5469,G5470,G5471,G5472,G5473,G5474,G5475,G5476,G5477,G5478,G5479,G5480,
       G5481,G5482,G5483,G5484,G5485,G5486,G5487,G5488,G5489,G5490,G5491,G5492,G5493,G5494,G5495,G5496,G5497,G5498,G5499,G5500,
       G5501,G5502,G5503,G5504,G5505,G5506,G5507,G5508,G5509,G5510,G5511,G5512,G5513,G5514,G5515,G5516,G5517,G5518,G5519,G5520,
       G5521,G5522,G5523,G5524,G5525,G5526,G5527,G5528,G5529,G5530,G5531,G5532,G5533,G5534,G5535,G5536,G5537,G5538,G5539,G5540,
       G5541,G5542,G5543,G5544,G5545,G5546,G5547,G5548,G5549,G5550,G5551,G5552,G5553,G5554,G5555,G5556,G5557,G5558,G5559,G5560,
       G5561,G5562,G5563,G5564,G5565,G5566,G5567,G5568,G5569,G5570,G5571,G5572,G5573,G5574,G5575,G5576,G5577,G5578,G5579,G5580,
       G5581,G5582,G5583,G5584,G5585,G5586,G5587,G5588,G5589,G5590,G5591,G5592,G5593,G5594,G5595,G5596,G5597,G5598,G5599,G5600,
       G5601,G5602,G5603,G5604,G5605,G5606,G5607,G5608,G5609,G5610,G5611,G5612,G5613,G5614,G5615,G5616,G5617,G5618,G5619,G5620,
       G5621,G5622,G5623,G5624,G5625,G5626,G5627,G5628,G5629,G5630,G5631,G5632,G5633,G5634,G5635,G5636,G5637,G5638,G5639,G5640,
       G5641,G5642,G5643,G5644,G5645,G5646,G5647,G5648,G5649,G5650,G5651,G5652,G5653,G5654,G5655,G5656,G5657,G5658,G5659,G5660,
       G5661,G5662,G5663,G5664,G5665,G5666,G5667,G5668,G5669,G5670,G5671,G5672,G5673,G5674,G5675,G5676,G5677,G5678,G5679,G5680,
       G5681,G5682,G5683,G5684,G5685,G5686,G5687,G5688,G5689,G5690,G5691,G5692,G5693,G5694,G5695,G5696,G5697,G5698,G5699,G5700,
       G5701,G5702,G5703,G5704,G5705,G5706,G5707,G5708,G5709,G5710,G5711,G5712,G5713,G5714,G5715,G5716,G5717,G5718,G5719,G5720,
       G5721,G5722,G5723,G5724,G5725,G5726,G5727,G5728,G5729,G5730,G5731,G5732,G5733,G5734,G5735,G5736,G5737,G5738,G5739,G5740,
       G5741,G5742,G5743,G5744,G5745,G5746,G5747,G5748,G5749,G5750,G5751,G5752,G5753,G5754,G5755,G5756,G5757,G5758,G5759,G5760,
       G5761,G5762,G5763,G5764,G5765,G5766,G5767,G5768,G5769,G5770,G5771,G5772,G5773,G5774,G5775,G5776,G5777,G5778,G5779,G5780,
       G5781,G5782,G5783,G5784,G5785,G5786,G5787,G5788,G5789,G5790,G5791,G5792,G5793,G5794,G5795,G5796,G5797,G5798,G5799,G5800,
       G5801,G5802,G5803,G5804,G5805,G5806,G5807,G5808,G5809,G5810,G5811,G5812,G5813,G5814,G5815,G5816,G5817,G5818,G5819,G5820,
       G5821,G5822,G5823,G5824,G5825,G5826,G5827,G5828,G5829,G5830,G5831,G5832,G5833,G5834,G5835,G5836,G5837,G5838,G5839,G5840,
       G5841,G5842,G5843,G5844,G5845,G5846,G5847,G5848,G5849,G5850,G5851,G5852,G5853,G5854,G5855,G5856,G5857,G5858,G5859,G5860,
       G5861,G5862,G5863,G5864,G5865,G5866,G5867,G5868,G5869,G5870,G5871,G5872,G5873,G5874,G5875,G5876,G5877,G5878,G5879,G5880,
       G5881,G5882,G5883,G5884,G5885,G5886,G5887,G5888,G5889,G5890,G5891,G5892,G5893,G5894,G5895,G5896,G5897,G5898,G5899,G5900,
       G5901,G5902,G5903,G5904,G5905,G5906,G5907,G5908,G5909,G5910,G5911,G5912,G5913,G5914,G5915,G5916,G5917,G5918,G5919,G5920,
       G5921,G5922,G5923,G5924,G5925,G5926,G5927,G5928,G5929,G5930,G5931,G5932,G5933,G5934,G5935,G5936,G5937,G5938,G5939,G5940,
       G5941,G5942,G5943,G5944,G5945,G5946,G5947,G5948,G5949,G5950,G5951,G5952,G5953,G5954,G5955,G5956,G5957,G5958,G5959,G5960,
       G5961,G5962,G5963,G5964,G5965,G5966,G5967,G5968,G5969,G5970,G5971,G5972,G5973,G5974,G5975,G5976,G5977,G5978,G5979,G5980,
       G5981,G5982,G5983,G5984,G5985,G5986,G5987,G5988,G5989,G5990,G5991,G5992,G5993,G5994,G5995,G5996,G5997,G5998,G5999,G6000,
       G6001,G6002,G6003,G6004,G6005,G6006,G6007,G6008,G6009,G6010,G6011,G6012,G6013,G6014,G6015,G6016,G6017,G6018,G6019,G6020,
       G6021,G6022,G6023,G6024,G6025,G6026,G6027,G6028,G6029,G6030,G6031,G6032,G6033,G6034,G6035,G6036,G6037,G6038,G6039,G6040,
       G6041,G6042,G6043,G6044,G6045,G6046,G6047,G6048,G6049,G6050,G6051,G6052,G6053,G6054,G6055,G6056,G6057,G6058,G6059,G6060,
       G6061,G6062,G6063,G6064,G6065,G6066,G6067,G6068,G6069,G6070,G6071,G6072,G6073,G6074,G6075,G6076,G6077,G6078,G6079,G6080,
       G6081,G6082,G6083,G6084,G6085,G6086,G6087,G6088,G6089,G6090,G6091,G6092,G6093,G6094,G6095,G6096,G6097,G6098,G6099,G6100,
       G6101,G6102,G6103,G6104,G6105,G6106,G6107,G6108,G6109,G6110,G6111,G6112,G6113,G6114,G6115,G6116,G6117,G6118,G6119,G6120,
       G6121,G6122,G6123,G6124,G6125,G6126,G6127,G6128,G6129,G6130,G6131,G6132,G6133,G6134,G6135,G6136,G6137,G6138,G6139,G6140,
       G6141,G6142,G6143,G6144,G6145,G6146,G6147,G6148,G6149,G6150,G6151,G6152,G6153,G6154,G6155,G6156,G6157,G6158,G6159,G6160,
       G6161,G6162,G6163,G6164,G6165,G6166,G6167,G6168,G6169,G6170,G6171,G6172,G6173,G6174,G6175,G6176,G6177,G6178,G6179,G6180,
       G6181,G6182,G6183,G6184,G6185,G6186,G6187,G6188,G6189,G6190,G6191,G6192,G6193,G6194,G6195,G6196,G6197,G6198,G6199,G6200,
       G6201,G6202,G6203,G6204,G6205,G6206,G6207,G6208,G6209,G6210,G6211,G6212,G6213,G6214,G6215,G6216,G6217,G6218,G6219,G6220,
       G6221,G6222,G6223,G6224,G6225,G6226,G6227,G6228,G6229,G6230,G6231,G6232,G6233,G6234,G6235,G6236,G6237,G6238,G6239,G6240,
       G6241,G6242,G6243,G6244,G6245,G6246,G6247,G6248,G6249,G6250,G6251,G6252,G6253,G6254,G6255,G6256,G6257,G6258,G6259,G6260,
       G6261,G6262,G6263,G6264,G6265,G6266,G6267,G6268,G6269,G6270,G6271,G6272,G6273,G6274,G6275,G6276,G6277,G6278,G6279,G6280,
       G6281,G6282,G6283,G6284,G6285,G6286,G6287,G6288,G6289,G6290,G6291,G6292,G6293,G6294,G6295,G6296,G6297,G6298,G6299,G6300,
       G6301,G6302,G6303,G6304,G6305,G6306,G6307,G6308,G6309,G6310,G6311,G6312,G6313,G6314,G6315,G6316,G6317,G6318,G6319,G6320,
       G6321,G6322,G6323,G6324,G6325,G6326,G6327,G6328,G6329,G6330,G6331,G6332,G6333,G6334,G6335,G6336,G6337,G6338,G6339,G6340,
       G6341,G6342,G6343,G6344,G6345,G6346,G6347,G6348,G6349,G6350,G6351,G6352,G6353,G6354,G6355,G6356,G6357,G6358,G6359,G6360,
       G6361,G6362,G6363,G6364,G6365,G6366,G6367,G6368,G6369,G6370,G6371,G6372,G6373,G6374,G6375,G6376,G6377,G6378,G6379,G6380,
       G6381,G6382,G6383,G6384,G6385,G6386,G6387,G6388,G6389,G6390,G6391,G6392,G6393,G6394,G6395,G6396,G6397,G6398,G6399,G6400,
       G6401,G6402,G6403,G6404,G6405,G6406,G6407,G6408,G6409,G6410,G6411,G6412,G6413,G6414,G6415,G6416,G6417,G6418,G6419,G6420,
       G6421,G6422,G6423,G6424,G6425,G6426,G6427,G6428,G6429,G6430,G6431,G6432,G6433,G6434,G6435,G6436,G6437,G6438,G6439,G6440,
       G6441,G6442,G6443,G6444,G6445,G6446,G6447,G6448,G6449,G6450,G6451,G6452,G6453,G6454,G6455,G6456,G6457,G6458,G6459,G6460,
       G6461,G6462,G6463,G6464,G6465,G6466,G6467,G6468,G6469,G6470,G6471,G6472,G6473,G6474,G6475,G6476,G6477,G6478,G6479,G6480,
       G6481,G6482,G6483,G6484,G6485,G6486,G6487,G6488,G6489,G6490,G6491,G6492,G6493,G6494,G6495,G6496,G6497,G6498,G6499,G6500,
       G6501,G6502,G6503,G6504,G6505,G6506,G6507,G6508,G6509,G6510,G6511,G6512,G6513,G6514,G6515,G6516,G6517,G6518,G6519,G6520,
       G6521,G6522,G6523,G6524,G6525,G6526,G6527,G6528,G6529,G6530,G6531,G6532,G6533,G6534,G6535,G6536,G6537,G6538,G6539,G6540,
       G6541,G6542,G6543,G6544,G6545,G6546,G6547,G6548,G6549,G6550,G6551,G6552,G6553,G6554,G6555,G6556,G6557,G6558,G6559,G6560,
       G6561,G6562,G6563,G6564,G6565,G6566,G6567,G6568,G6569,G6570,G6571,G6572,G6573,G6574,G6575,G6576,G6577,G6578,G6579,G6580,
       G6581,G6582,G6583,G6584,G6585,G6586,G6587,G6588,G6589,G6590,G6591,G6592,G6593,G6594,G6595,G6596,G6597,G6598,G6599,G6600,
       G6601,G6602,G6603,G6604,G6605,G6606,G6607,G6608,G6609,G6610,G6611,G6612,G6613,G6614,G6615,G6616,G6617,G6618,G6619,G6620,
       G6621,G6622,G6623,G6624,G6625,G6626,G6627,G6628,G6629,G6630,G6631,G6632,G6633,G6634,G6635,G6636,G6637,G6638,G6639,G6640,
       G6641,G6642,G6643,G6644,G6645,G6646,G6647,G6648,G6649,G6650,G6651,G6652,G6653,G6654,G6655,G6656,G6657,G6658,G6659,G6660,
       G6661,G6662,G6663,G6664,G6665,G6666,G6667,G6668,G6669,G6670,G6671,G6672,G6673,G6674,G6675,G6676,G6677,G6678,G6679,G6680,
       G6681,G6682,G6683,G6684,G6685,G6686,G6687,G6688,G6689,G6690,G6691,G6692,G6693,G6694,G6695,G6696,G6697,G6698,G6699,G6700,
       G6701,G6702,G6703,G6704,G6705,G6706,G6707,G6708,G6709,G6710,G6711,G6712,G6713,G6714,G6715,G6716,G6717,G6718,G6719,G6720,
       G6721,G6722,G6723,G6724,G6725,G6726,G6727,G6728,G6729,G6730,G6731,G6732,G6733,G6734,G6735,G6736,G6737,G6738,G6739,G6740,
       G6741,G6742,G6743,G6744,G6745,G6746,G6747,G6748,G6749,G6750,G6751,G6752,G6753,G6754,G6755,G6756,G6757,G6758,G6759,G6760,
       G6761,G6762,G6763,G6764,G6765,G6766,G6767,G6768,G6769,G6770,G6771,G6772,G6773,G6774,G6775,G6776,G6777,G6778,G6779,G6780,
       G6781,G6782,G6783,G6784,G6785,G6786,G6787,G6788,G6789,G6790,G6791,G6792,G6793,G6794,G6795,G6796,G6797,G6798,G6799,G6800,
       G6801,G6802,G6803,G6804,G6805,G6806,G6807,G6808,G6809,G6810,G6811,G6812,G6813,G6814,G6815,G6816,G6817,G6818,G6819,G6820,
       G6821,G6822,G6823,G6824,G6825,G6826,G6827,G6828,G6829,G6830,G6831,G6832,G6833,G6834,G6835,G6836,G6837,G6838,G6839,G6840,
       G6841,G6842,G6843,G6844,G6845,G6846,G6847,G6848,G6849,G6850,G6851,G6852,G6853,G6854,G6855,G6856,G6857,G6858,G6859,G6860,
       G6861,G6862,G6863,G6864,G6865,G6866,G6867,G6868,G6869,G6870,G6871,G6872,G6873,G6874,G6875,G6876,G6877,G6878,G6879,G6880,
       G6881,G6882,G6883,G6884,G6885,G6886,G6887,G6888,G6889,G6890,G6891,G6892,G6893,G6894,G6895,G6896,G6897,G6898,G6899,G6900,
       G6901,G6902,G6903,G6904,G6905,G6906,G6907,G6908,G6909,G6910,G6911,G6912,G6913,G6914,G6915,G6916,G6917,G6918,G6919,G6920,
       G6921,G6922,G6923,G6924,G6925,G6926,G6927,G6928,G6929,G6930,G6931,G6932,G6933,G6934,G6935,G6936,G6937,G6938,G6939,G6940,
       G6941,G6942,G6943,G6944,G6945,G6946,G6947,G6948,G6949,G6950,G6951,G6952,G6953,G6954,G6955,G6956,G6957,G6958,G6959,G6960,
       G6961,G6962,G6963,G6964,G6965,G6966,G6967,G6968,G6969,G6970,G6971,G6972,G6973,G6974,G6975,G6976,G6977,G6978,G6979,G6980,
       G6981,G6982,G6983,G6984,G6985,G6986,G6987,G6988,G6989,G6990,G6991,G6992,G6993,G6994,G6995,G6996,G6997,G6998,G6999,G7000,
       G7001,G7002,G7003,G7004,G7005,G7006,G7007,G7008,G7009,G7010,G7011,G7012,G7013,G7014,G7015,G7016,G7017,G7018,G7019,G7020,
       G7021,G7022,G7023,G7024,G7025,G7026,G7027,G7028,G7029,G7030,G7031,G7032,G7033,G7034,G7035,G7036,G7037,G7038,G7039,G7040,
       G7041,G7042,G7043,G7044,G7045,G7046,G7047,G7048,G7049,G7050,G7051,G7052,G7053,G7054,G7055,G7056,G7057,G7058,G7059,G7060,
       G7061,G7062,G7063,G7064,G7065,G7066,G7067,G7068,G7069,G7070,G7071,G7072,G7073,G7074,G7075,G7076,G7077,G7078,G7079,G7080,
       G7081,G7082,G7083,G7084,G7085,G7086,G7087,G7088,G7089,G7090,G7091,G7092,G7093,G7094,G7095,G7096,G7097,G7098,G7099,G7100,
       G7101,G7102,G7103,G7104,G7105,G7106,G7107,G7108,G7109,G7110,G7111,G7112,G7113,G7114,G7115,G7116,G7117,G7118,G7119,G7120,
       G7121,G7122,G7123,G7124,G7125,G7126,G7127,G7128,G7129,G7130,G7131,G7132,G7133,G7134,G7135,G7136,G7137,G7138,G7139,G7140,
       G7141,G7142,G7143,G7144,G7145,G7146,G7147,G7148,G7149,G7150,G7151,G7152,G7153,G7154,G7155,G7156,G7157,G7158,G7159,G7160,
       G7161,G7162,G7163,G7164,G7165,G7166,G7167,G7168,G7169,G7170,G7171,G7172,G7173,G7174,G7175,G7176,G7177,G7178,G7179,G7180,
       G7181,G7182,G7183,G7184,G7185,G7186,G7187,G7188,G7189,G7190,G7191,G7192,G7193,G7194,G7195,G7196,G7197,G7198,G7199,G7200,
       G7201,G7202,G7203,G7204,G7205,G7206,G7207,G7208,G7209,G7210,G7211,G7212,G7213,G7214,G7215,G7216,G7217,G7218,G7219,G7220,
       G7221,G7222,G7223,G7224,G7225,G7226,G7227,G7228,G7229,G7230,G7231,G7232,G7233,G7234,G7235,G7236,G7237,G7238,G7239,G7240,
       G7241,G7242,G7243,G7244,G7245,G7246,G7247,G7248,G7249,G7250,G7251,G7252,G7253,G7254,G7255,G7256,G7257,G7258,G7259,G7260,
       G7261,G7262,G7263,G7264,G7265,G7266,G7267,G7268,G7269,G7270,G7271,G7272,G7273,G7274,G7275,G7276,G7277,G7278,G7279,G7280,
       G7281,G7282,G7283,G7284,G7285,G7286,G7287,G7288,G7289,G7290,G7291,G7292,G7293,G7294,G7295,G7296,G7297,G7298,G7299,G7300,
       G7301,G7302,G7303,G7304,G7305,G7306,G7307,G7308,G7309,G7310,G7311,G7312,G7313,G7314,G7315,G7316,G7317,G7318,G7319,G7320,
       G7321,G7322,G7323,G7324,G7325,G7326,G7327,G7328,G7329,G7330,G7331,G7332,G7333,G7334,G7335,G7336,G7337,G7338,G7339,G7340,
       G7341,G7342,G7343,G7344,G7345,G7346,G7347,G7348,G7349,G7350,G7351,G7352,G7353,G7354,G7355,G7356,G7357,G7358,G7359,G7360,
       G7361,G7362,G7363,G7364,G7365,G7366,G7367,G7368,G7369,G7370,G7371,G7372,G7373,G7374,G7375,G7376,G7377,G7378,G7379,G7380,
       G7381,G7382,G7383,G7384,G7385,G7386,G7387,G7388,G7389,G7390,G7391,G7392,G7393,G7394,G7395,G7396,G7397,G7398,G7399,G7400,
       G7401,G7402,G7403,G7404,G7405,G7406,G7407,G7408,G7409,G7410,G7411,G7412,G7413,G7414,G7415,G7416,G7417,G7418,G7419,G7420,
       G7421,G7422,G7423,G7424,G7425,G7426,G7427,G7428,G7429,G7430,G7431,G7432,G7433,G7434,G7435,G7436,G7437,G7438,G7439,G7440,
       G7441,G7442,G7443,G7444,G7445,G7446,G7447,G7448,G7449,G7450,G7451,G7452,G7453,G7454,G7455,G7456,G7457,G7458,G7459,G7460,
       G7461,G7462,G7463,G7464,G7465,G7466,G7467,G7468,G7469,G7470,G7471,G7472,G7473,G7474,G7475,G7476,G7477,G7478,G7479,G7480,
       G7481,G7482,G7483,G7484,G7485,G7486,G7487,G7488,G7489,G7490,G7491,G7492,G7493,G7494,G7495,G7496,G7497,G7498,G7499,G7500,
       G7501,G7502,G7503,G7504,G7505,G7506,G7507,G7508,G7509,G7510,G7511,G7512,G7513,G7514,G7515,G7516,G7517,G7518,G7519,G7520,
       G7521,G7522,G7523,G7524,G7525,G7526,G7527,G7528,G7529,G7530,G7531,G7532,G7533,G7534,G7535,G7536,G7537,G7538,G7539,G7540,
       G7541,G7542,G7543,G7544,G7545,G7546,G7547,G7548,G7549,G7550,G7551,G7552,G7553,G7554,G7555,G7556,G7557,G7558,G7559,G7560,
       G7561,G7562,G7563,G7564,G7565,G7566,G7567,G7568,G7569,G7570,G7571,G7572,G7573,G7574,G7575,G7576,G7577,G7578,G7579,G7580,
       G7581,G7582,G7583,G7584,G7585,G7586,G7587,G7588,G7589,G7590,G7591,G7592,G7593,G7594,G7595,G7596,G7597,G7598,G7599,G7600,
       G7601,G7602,G7603,G7604,G7605,G7606,G7607,G7608,G7609,G7610,G7611,G7612,G7613,G7614,G7615,G7616,G7617,G7618,G7619,G7620,
       G7621,G7622,G7623,G7624,G7625,G7626,G7627,G7628,G7629,G7630,G7631,G7632,G7633,G7634,G7635,G7636,G7637,G7638,G7639,G7640,
       G7641,G7642,G7643,G7644,G7645,G7646,G7647,G7648,G7649,G7650,G7651,G7652,G7653,G7654,G7655,G7656,G7657,G7658,G7659,G7660,
       G7661,G7662,G7663,G7664,G7665,G7666,G7667,G7668,G7669,G7670,G7671,G7672,G7673,G7674,G7675,G7676,G7677,G7678,G7679,G7680,
       G7681,G7682,G7683,G7684,G7685,G7686,G7687,G7688,G7689,G7690,G7691,G7692,G7693,G7694,G7695,G7696,G7697,G7698,G7699,G7700,
       G7701,G7702,G7703,G7704,G7705,G7706,G7707,G7708,G7709,G7710,G7711,G7712,G7713,G7714,G7715,G7716,G7717,G7718,G7719,G7720,
       G7721,G7722,G7723,G7724,G7725,G7726,G7727,G7728,G7729,G7730,G7731,G7732,G7733,G7734,G7735,G7736,G7737,G7738,G7739,G7740,
       G7741,G7742,G7743,G7744,G7745,G7746,G7747,G7748,G7749,G7750,G7751,G7752,G7753,G7754,G7755,G7756,G7757,G7758,G7759,G7760,
       G7761,G7762,G7763,G7764,G7765,G7766,G7767,G7768,G7769,G7770,G7771,G7772,G7773,G7774,G7775,G7776,G7777,G7778,G7779,G7780,
       G7781,G7782,G7783,G7784,G7785,G7786,G7787,G7788,G7789,G7790,G7791,G7792,G7793,G7794,G7795,G7796,G7797,G7798,G7799,G7800,
       G7801,G7802,G7803,G7804,G7805,G7806,G7807,G7808,G7809,G7810,G7811,G7812,G7813,G7814,G7815,G7816,G7817,G7818,G7819,G7820,
       G7821,G7822,G7823,G7824,G7825,G7826,G7827,G7828,G7829,G7830,G7831,G7832,G7833,G7834,G7835,G7836,G7837,G7838,G7839,G7840,
       G7841,G7842,G7843,G7844,G7845,G7846,G7847,G7848,G7849,G7850,G7851,G7852,G7853,G7854,G7855,G7856,G7857,G7858,G7859,G7860,
       G7861,G7862,G7863,G7864,G7865,G7866,G7867,G7868,G7869,G7870,G7871,G7872,G7873,G7874,G7875,G7876,G7877,G7878,G7879,G7880,
       G7881,G7882,G7883,G7884,G7885,G7886,G7887,G7888,G7889,G7890,G7891,G7892,G7893,G7894,G7895,G7896,G7897,G7898,G7899,G7900,
       G7901,G7902,G7903,G7904,G7905,G7906,G7907,G7908,G7909,G7910,G7911,G7912,G7913,G7914,G7915,G7916,G7917,G7918,G7919,G7920,
       G7921,G7922,G7923,G7924,G7925,G7926,G7927,G7928,G7929,G7930,G7931,G7932,G7933,G7934,G7935,G7936,G7937,G7938,G7939,G7940,
       G7941,G7942,G7943,G7944,G7945,G7946,G7947,G7948,G7949,G7950,G7951,G7952,G7953,G7954,G7955,G7956,G7957,G7958,G7959,G7960,
       G7961,G7962,G7963,G7964,G7965,G7966,G7967,G7968,G7969,G7970,G7971,G7972,G7973,G7974,G7975,G7976,G7977,G7978,G7979,G7980,
       G7981,G7982,G7983,G7984,G7985,G7986,G7987,G7988,G7989,G7990,G7991,G7992,G7993,G7994,G7995,G7996,G7997,G7998,G7999,G8000,
       G8001,G8002,G8003,G8004,G8005,G8006,G8007,G8008,G8009,G8010,G8011,G8012,G8013,G8014,G8015,G8016,G8017,G8018,G8019,G8020,
       G8021,G8022,G8023,G8024,G8025,G8026,G8027,G8028,G8029,G8030,G8031,G8032,G8033,G8034,G8035,G8036,G8037,G8038,G8039,G8040,
       G8041,G8042,G8043,G8044,G8045,G8046,G8047,G8048,G8049,G8050,G8051,G8052,G8053,G8054,G8055,G8056,G8057,G8058,G8059,G8060,
       G8061,G8062,G8063,G8064,G8065,G8066,G8067,G8068,G8069,G8070,G8071,G8072,G8073,G8074,G8075,G8076,G8077,G8078,G8079,G8080,
       G8081,G8082,G8083,G8084,G8085,G8086,G8087,G8088,G8089,G8090,G8091,G8092,G8093,G8094,G8095,G8096,G8097,G8098,G8099,G8100,
       G8101,G8102,G8103,G8104,G8105,G8106,G8107,G8108,G8109,G8110,G8111,G8112,G8113,G8114,G8115,G8116,G8117,G8118,G8119,G8120,
       G8121,G8122,G8123,G8124,G8125,G8126,G8127,G8128,G8129,G8130,G8131,G8132,G8133,G8134,G8135,G8136,G8137,G8138,G8139,G8140,
       G8141,G8142,G8143,G8144,G8145,G8146,G8147,G8148,G8149,G8150,G8151,G8152,G8153,G8154,G8155,G8156,G8157,G8158,G8159,G8160,
       G8161,G8162,G8163,G8164,G8165,G8166,G8167,G8168,G8169,G8170,G8171,G8172,G8173,G8174,G8175,G8176,G8177,G8178,G8179,G8180,
       G8181,G8182,G8183,G8184,G8185,G8186,G8187,G8188,G8189,G8190,G8191,G8192,G8193,G8194,G8195,G8196,G8197,G8198,G8199,G8200,
       G8201,G8202,G8203,G8204,G8205,G8206,G8207,G8208,G8209,G8210,G8211,G8212,G8213,G8214,G8215,G8216,G8217,G8218,G8219,G8220,
       G8221,G8222,G8223,G8224,G8225,G8226,G8227,G8228,G8229,G8230,G8231,G8232,G8233,G8234,G8235,G8236,G8237,G8238,G8239,G8240,
       G8241,G8242,G8243,G8244,G8245,G8246,G8247,G8248,G8249,G8250,G8251,G8252,G8253,G8254,G8255,G8256,G8257,G8258,G8259,G8260,
       G8261,G8262,G8263,G8264,G8265,G8266,G8267,G8268,G8269,G8270,G8271,G8272,G8273,G8274,G8275,G8276,G8277,G8278,G8279,G8280,
       G8281,G8282,G8283,G8284,G8285,G8286,G8287,G8288,G8289,G8290,G8291,G8292,G8293,G8294,G8295,G8296,G8297,G8298,G8299,G8300,
       G8301,G8302,G8303,G8304,G8305,G8306,G8307,G8308,G8309,G8310,G8311,G8312,G8313,G8314,G8315,G8316,G8317,G8318,G8319,G8320,
       G8321,G8322,G8323,G8324,G8325,G8326,G8327,G8328,G8329,G8330,G8331,G8332,G8333,G8334,G8335,G8336,G8337,G8338,G8339,G8340,
       G8341,G8342,G8343,G8344,G8345,G8346,G8347,G8348,G8349,G8350,G8351,G8352,G8353,G8354,G8355,G8356,G8357,G8358,G8359,G8360,
       G8361,G8362,G8363,G8364,G8365,G8366,G8367,G8368,G8369,G8370,G8371,G8372,G8373,G8374,G8375,G8376,G8377,G8378,G8379,G8380,
       G8381,G8382,G8383,G8384,G8385,G8386,G8387,G8388,G8389,G8390,G8391,G8392,G8393,G8394,G8395,G8396,G8397,G8398,G8399,G8400,
       G8401,G8402,G8403,G8404,G8405,G8406,G8407,G8408,G8409,G8410,G8411,G8412,G8413,G8414,G8415,G8416,G8417,G8418,G8419,G8420,
       G8421,G8422,G8423,G8424,G8425,G8426,G8427,G8428,G8429,G8430,G8431,G8432,G8433,G8434,G8435,G8436,G8437,G8438,G8439,G8440,
       G8441,G8442,G8443,G8444,G8445,G8446,G8447,G8448,G8449,G8450,G8451,G8452,G8453,G8454,G8455,G8456,G8457,G8458,G8459,G8460,
       G8461,G8462,G8463,G8464,G8465,G8466,G8467,G8468,G8469,G8470,G8471,G8472,G8473,G8474,G8475,G8476,G8477,G8478,G8479,G8480,
       G8481,G8482,G8483,G8484,G8485,G8486,G8487,G8488,G8489,G8490,G8491,G8492,G8493,G8494,G8495,G8496,G8497,G8498,G8499,G8500,
       G8501,G8502,G8503,G8504,G8505,G8506,G8507,G8508,G8509,G8510,G8511,G8512,G8513,G8514,G8515,G8516,G8517,G8518,G8519,G8520,
       G8521,G8522,G8523,G8524,G8525,G8526,G8527,G8528,G8529,G8530,G8531,G8532,G8533,G8534,G8535,G8536,G8537,G8538,G8539,G8540,
       G8541,G8542,G8543,G8544,G8545,G8546,G8547,G8548,G8549,G8550,G8551,G8552,G8553,G8554,G8555,G8556,G8557,G8558,G8559,G8560,
       G8561,G8562,G8563,G8564,G8565,G8566,G8567,G8568,G8569,G8570,G8571,G8572,G8573,G8574,G8575,G8576,G8577,G8578,G8579,G8580,
       G8581,G8582,G8583,G8584,G8585,G8586,G8587,G8588,G8589,G8590,G8591,G8592,G8593,G8594,G8595,G8596,G8597,G8598,G8599,G8600,
       G8601,G8602,G8603,G8604,G8605,G8606,G8607,G8608,G8609,G8610,G8611,G8612,G8613,G8614,G8615,G8616,G8617,G8618,G8619,G8620,
       G8621,G8622,G8623,G8624,G8625,G8626,G8627,G8628,G8629,G8630,G8631,G8632,G8633,G8634,G8635,G8636,G8637,G8638,G8639,G8640,
       G8641,G8642,G8643,G8644,G8645,G8646,G8647,G8648,G8649,G8650,G8651,G8652,G8653,G8654,G8655,G8656,G8657,G8658,G8659,G8660,
       G8661,G8662,G8663,G8664,G8665,G8666,G8667,G8668,G8669,G8670,G8671,G8672,G8673,G8674,G8675,G8676,G8677,G8678,G8679,G8680,
       G8681,G8682,G8683,G8684,G8685,G8686,G8687,G8688,G8689,G8690,G8691,G8692,G8693,G8694,G8695,G8696,G8697,G8698,G8699,G8700,
       G8701,G8702,G8703,G8704,G8705,G8706,G8707,G8708,G8709,G8710,G8711,G8712,G8713,G8714,G8715,G8716,G8717,G8718,G8719,G8720,
       G8721,G8722,G8723,G8724,G8725,G8726,G8727,G8728,G8729,G8730,G8731,G8732,G8733,G8734,G8735,G8736,G8737,G8738,G8739,G8740,
       G8741,G8742,G8743,G8744,G8745,G8746,G8747,G8748,G8749,G8750,G8751,G8752,G8753,G8754,G8755,G8756,G8757,G8758,G8759,G8760,
       G8761,G8762,G8763,G8764,G8765,G8766,G8767,G8768,G8769,G8770,G8771,G8772,G8773,G8774,G8775,G8776,G8777,G8778,G8779,G8780,
       G8781,G8782,G8783,G8784,G8785,G8786,G8787,G8788,G8789,G8790,G8791,G8792,G8793,G8794,G8795,G8796,G8797,G8798,G8799,G8800,
       G8801,G8802,G8803,G8804,G8805,G8806,G8807,G8808,G8809,G8810,G8811,G8812,G8813,G8814,G8815,G8816,G8817,G8818,G8819,G8820,
       G8821,G8822,G8823,G8824,G8825,G8826,G8827,G8828,G8829,G8830,G8831,G8832,G8833,G8834,G8835,G8836,G8837,G8838,G8839,G8840,
       G8841,G8842,G8843,G8844,G8845,G8846,G8847,G8848,G8849,G8850,G8851,G8852,G8853,G8854,G8855,G8856,G8857,G8858,G8859,G8860,
       G8861,G8862,G8863,G8864,G8865,G8866,G8867,G8868,G8869,G8870,G8871,G8872,G8873,G8874,G8875,G8876,G8877,G8878,G8879,G8880,
       G8881,G8882,G8883,G8884,G8885,G8886,G8887,G8888,G8889,G8890,G8891,G8892,G8893,G8894,G8895,G8896,G8897,G8898,G8899,G8900,
       G8901,G8902,G8903,G8904,G8905,G8906,G8907,G8908,G8909,G8910,G8911,G8912,G8913,G8914,G8915,G8916,G8917,G8918,G8919,G8920,
       G8921,G8922,G8923,G8924,G8925,G8926,G8927,G8928,G8929,G8930,G8931,G8932,G8933,G8934,G8935,G8936,G8937,G8938,G8939,G8940,
       G8941,G8942,G8943,G8944,G8945,G8946,G8947,G8948,G8949,G8950,G8951,G8952,G8953,G8954,G8955,G8956,G8957,G8958,G8959,G8960,
       G8961,G8962,G8963,G8964,G8965,G8966,G8967,G8968,G8969,G8970,G8971,G8972,G8973,G8974,G8975,G8976,G8977,G8978,G8979,G8980,
       G8981,G8982,G8983,G8984,G8985,G8986,G8987,G8988,G8989,G8990,G8991,G8992,G8993,G8994,G8995,G8996,G8997,G8998,G8999,G9000,
       G9001,G9002,G9003,G9004,G9005,G9006,G9007,G9008,G9009,G9010,G9011,G9012,G9013,G9014,G9015,G9016,G9017,G9018,G9019,G9020,
       G9021,G9022,G9023,G9024,G9025,G9026,G9027,G9028,G9029,G9030,G9031,G9032,G9033,G9034,G9035,G9036,G9037,G9038,G9039,G9040,
       G9041,G9042,G9043,G9044,G9045,G9046,G9047,G9048,G9049,G9050,G9051,G9052,G9053,G9054,G9055,G9056,G9057,G9058,G9059,G9060,
       G9061,G9062,G9063,G9064,G9065,G9066,G9067,G9068,G9069,G9070,G9071,G9072,G9073,G9074,G9075,G9076,G9077,G9078,G9079,G9080,
       G9081,G9082,G9083,G9084,G9085,G9086,G9087,G9088,G9089,G9090,G9091,G9092,G9093,G9094,G9095,G9096,G9097,G9098,G9099,G9100,
       G9101,G9102,G9103,G9104,G9105,G9106,G9107,G9108,G9109,G9110,G9111,G9112,G9113,G9114,G9115,G9116,G9117,G9118,G9119,G9120,
       G9121,G9122,G9123,G9124,G9125,G9126,G9127,G9128,G9129,G9130,G9131,G9132,G9133,G9134,G9135,G9136,G9137,G9138,G9139,G9140,
       G9141,G9142,G9143,G9144,G9145,G9146,G9147,G9148,G9149,G9150,G9151,G9152,G9153,G9154,G9155,G9156,G9157,G9158,G9159,G9160,
       G9161,G9162,G9163,G9164,G9165,G9166,G9167,G9168,G9169,G9170,G9171,G9172,G9173,G9174,G9175,G9176,G9177,G9178,G9179,G9180,
       G9181,G9182,G9183,G9184,G9185,G9186,G9187,G9188,G9189,G9190,G9191,G9192,G9193,G9194,G9195,G9196,G9197,G9198,G9199,G9200,
       G9201,G9202,G9203,G9204,G9205,G9206,G9207,G9208,G9209,G9210,G9211,G9212,G9213,G9214,G9215,G9216,G9217,G9218,G9219,G9220,
       G9221,G9222,G9223,G9224,G9225,G9226,G9227,G9228,G9229,G9230,G9231,G9232,G9233,G9234,G9235,G9236,G9237,G9238,G9239,G9240,
       G9241,G9242,G9243,G9244,G9245,G9246,G9247,G9248,G9249,G9250,G9251,G9252,G9253,G9254,G9255,G9256,G9257,G9258,G9259,G9260,
       G9261,G9262,G9263,G9264,G9265,G9266,G9267,G9268,G9269,G9270,G9271,G9272,G9273,G9274,G9275,G9276,G9277,G9278,G9279,G9280,
       G9281,G9282,G9283,G9284,G9285,G9286,G9287,G9288,G9289,G9290,G9291,G9292,G9293,G9294,G9295,G9296,G9297,G9298,G9299,G9300,
       G9301,G9302,G9303,G9304,G9305,G9306,G9307,G9308,G9309,G9310,G9311,G9312,G9313,G9314,G9315,G9316,G9317,G9318,G9319,G9320,
       G9321,G9322,G9323,G9324,G9325,G9326,G9327,G9328,G9329,G9330,G9331,G9332,G9333,G9334,G9335,G9336,G9337,G9338,G9339,G9340,
       G9341,G9342,G9343,G9344,G9345,G9346,G9347,G9348,G9349,G9350,G9351,G9352,G9353,G9354,G9355,G9356,G9357,G9358,G9359,G9360,
       G9361,G9362,G9363,G9364,G9365,G9366,G9367,G9368,G9369,G9370,G9371,G9372,G9373,G9374,G9375,G9376,G9377,G9378,G9379,G9380,
       G9381,G9382,G9383,G9384,G9385,G9386,G9387,G9388,G9389,G9390,G9391,G9392,G9393,G9394,G9395,G9396,G9397,G9398,G9399,G9400,
       G9401,G9402,G9403,G9404,G9405,G9406,G9407,G9408,G9409,G9410,G9411,G9412,G9413,G9414,G9415,G9416,G9417,G9418,G9419,G9420,
       G9421,G9422,G9423,G9424,G9425,G9426,G9427,G9428,G9429,G9430,G9431,G9432,G9433,G9434,G9435,G9436,G9437,G9438,G9439,G9440,
       G9441,G9442,G9443,G9444,G9445,G9446,G9447,G9448,G9449,G9450,G9451,G9452,G9453,G9454,G9455,G9456,G9457,G9458,G9459,G9460,
       G9461,G9462,G9463,G9464,G9465,G9466,G9467,G9468,G9469,G9470,G9471,G9472,G9473,G9474,G9475,G9476,G9477,G9478,G9479,G9480,
       G9481,G9482,G9483,G9484,G9485,G9486,G9487,G9488,G9489,G9490,G9491,G9492,G9493,G9494,G9495,G9496,G9497,G9498,G9499,G9500,
       G9501,G9502,G9503,G9504,G9505,G9506,G9507,G9508,G9509,G9510,G9511,G9512,G9513,G9514,G9515,G9516,G9517,G9518,G9519,G9520,
       G9521,G9522,G9523,G9524,G9525,G9526,G9527,G9528,G9529,G9530,G9531,G9532,G9533,G9534,G9535,G9536,G9537,G9538,G9539,G9540,
       G9541,G9542,G9543,G9544,G9545,G9546,G9547,G9548,G9549,G9550,G9551,G9552,G9553,G9554,G9555,G9556,G9557,G9558,G9559,G9560,
       G9561,G9562,G9563,G9564,G9565,G9566,G9567,G9568,G9569,G9570,G9571,G9572,G9573,G9574,G9575,G9576,G9577,G9578,G9579,G9580,
       G9581,G9582,G9583,G9584,G9585,G9586,G9587,G9588,G9589,G9590,G9591,G9592,G9593,G9594,G9595,G9596,G9597,G9598,G9599,G9600,
       G9601,G9602,G9603,G9604,G9605,G9606,G9607,G9608,G9609,G9610,G9611,G9612,G9613,G9614,G9615,G9616,G9617,G9618,G9619,G9620,
       G9621,G9622,G9623,G9624,G9625,G9626,G9627,G9628,G9629,G9630,G9631,G9632,G9633,G9634,G9635,G9636,G9637,G9638,G9639,G9640,
       G9641,G9642,G9643,G9644,G9645,G9646,G9647,G9648,G9649,G9650,G9651,G9652,G9653,G9654,G9655,G9656,G9657,G9658,G9659,G9660,
       G9661,G9662,G9663,G9664,G9665,G9666,G9667,G9668,G9669,G9670,G9671,G9672,G9673,G9674,G9675,G9676,G9677,G9678,G9679,G9680,
       G9681,G9682,G9683,G9684,G9685,G9686,G9687,G9688,G9689,G9690,G9691,G9692,G9693,G9694,G9695,G9696,G9697,G9698,G9699,G9700,
       G9701,G9702,G9703,G9704,G9705,G9706,G9707,G9708,G9709,G9710,G9711,G9712,G9713,G9714,G9715,G9716,G9717,G9718,G9719,G9720,
       G9721,G9722,G9723,G9724,G9725,G9726,G9727,G9728,G9729,G9730,G9731,G9732,G9733,G9734,G9735,G9736,G9737,G9738,G9739,G9740,
       G9741,G9742,G9743,G9744,G9745,G9746,G9747,G9748,G9749,G9750,G9751,G9752,G9753,G9754,G9755,G9756,G9757,G9758,G9759,G9760,
       G9761,G9762,G9763,G9764,G9765,G9766,G9767,G9768,G9769,G9770,G9771,G9772,G9773,G9774,G9775,G9776,G9777,G9778,G9779,G9780,
       G9781,G9782,G9783,G9784,G9785,G9786,G9787,G9788,G9789,G9790,G9791,G9792,G9793,G9794,G9795,G9796,G9797,G9798,G9799,G9800,
       G9801,G9802,G9803,G9804,G9805,G9806,G9807,G9808,G9809,G9810,G9811,G9812,G9813,G9814,G9815,G9816,G9817,G9818,G9819,G9820,
       G9821,G9822,G9823,G9824,G9825,G9826,G9827,G9828,G9829,G9830,G9831,G9832,G9833,G9834,G9835,G9836,G9837,G9838,G9839,G9840,
       G9841,G9842,G9843,G9844,G9845,G9846,G9847,G9848,G9849,G9850,G9851,G9852,G9853,G9854,G9855,G9856,G9857,G9858,G9859,G9860,
       G9861,G9862,G9863,G9864,G9865,G9866,G9867,G9868,G9869,G9870,G9871,G9872,G9873,G9874,G9875,G9876,G9877,G9878,G9879,G9880,
       G9881,G9882,G9883,G9884,G9885,G9886,G9887,G9888,G9889,G9890,G9891,G9892,G9893,G9894,G9895,G9896,G9897,G9898,G9899,G9900,
       G9901,G9902,G9903,G9904,G9905,G9906,G9907,G9908,G9909,G9910,G9911,G9912,G9913,G9914,G9915,G9916,G9917,G9918,G9919,G9920,
       G9921,G9922,G9923,G9924,G9925,G9926,G9927,G9928,G9929,G9930,G9931,G9932,G9933,G9934,G9935,G9936,G9937,G9938,G9939,G9940,
       G9941,G9942,G9943,G9944,G9945,G9946,G9947,G9948,G9949,G9950,G9951,G9952,G9953,G9954,G9955,G9956,G9957,G9958,G9959,G9960,
       G9961,G9962,G9963,G9964,G9965,G9966,G9967,G9968,G9969,G9970,G9971,G9972,G9973,G9974,G9975,G9976,G9977,G9978,G9979,G9980,
       G9981,G9982,G9983,G9984,G9985,G9986,G9987,G9988,G9989,G9990,G9991,G9992,G9993,G9994,G9995,G9996,G9997,G9998,G9999,G10000,
       G10001,G10002,G10003,G10004,G10005,G10006,G10007,G10008,G10009,G10010,G10011,G10012,G10013,G10014,G10015,G10016,G10017,G10018,G10019,G10020,
       G10021,G10022,G10023,G10024,G10025,G10026,G10027,G10028,G10029,G10030,G10031,G10032,G10033,G10034,G10035,G10036,G10037,G10038,G10039,G10040,
       G10041,G10042,G10043,G10044,G10045,G10046,G10047,G10048,G10049,G10050,G10051,G10052,G10053,G10054,G10055,G10056,G10057,G10058,G10059,G10060,
       G10061,G10062,G10063,G10064,G10065,G10066,G10067,G10068,G10069,G10070,G10071,G10072,G10073,G10074,G10075,G10076,G10077,G10078,G10079,G10080,
       G10081,G10082,G10083,G10084,G10085,G10086,G10087,G10088,G10089,G10090,G10091,G10092,G10093,G10094,G10095,G10096,G10097,G10098,G10099,G10100,
       G10101,G10102,G10103,G10104,G10105,G10106,G10107,G10108,G10109,G10110,G10111,G10112,G10113,G10114,G10115,G10116,G10117,G10118,G10119,G10120,
       G10121,G10122,G10123,G10124,G10125,G10126,G10127,G10128,G10129,G10130,G10131,G10132,G10133,G10134,G10135,G10136,G10137,G10138,G10139,G10140,
       G10141,G10142,G10143,G10144,G10145,G10146,G10147,G10148,G10149,G10150,G10151,G10152,G10153,G10154,G10155,G10156,G10157,G10158,G10159,G10160,
       G10161,G10162,G10163,G10164,G10165,G10166,G10167,G10168,G10169,G10170,G10171,G10172,G10173,G10174,G10175,G10176,G10177,G10178,G10179,G10180,
       G10181,G10182,G10183,G10184,G10185,G10186,G10187,G10188,G10189,G10190,G10191,G10192,G10193,G10194,G10195,G10196,G10197,G10198,G10199,G10200,
       G10201,G10202,G10203,G10204,G10205,G10206,G10207,G10208,G10209,G10210,G10211,G10212,G10213,G10214,G10215,G10216,G10217,G10218,G10219,G10220,
       G10221,G10222,G10223,G10224,G10225,G10226,G10227,G10228,G10229,G10230,G10231,G10232,G10233,G10234,G10235,G10236,G10237,G10238,G10239,G10240,
       G10241,G10242,G10243,G10244,G10245,G10246,G10247,G10248,G10249,G10250,G10251,G10252,G10253,G10254,G10255,G10256,G10257,G10258,G10259,G10260,
       G10261,G10262,G10263,G10264,G10265,G10266,G10267,G10268,G10269,G10270,G10271,G10272,G10273,G10274,G10275,G10276,G10277,G10278,G10279,G10280,
       G10281,G10282,G10283,G10284,G10285,G10286,G10287,G10288,G10289,G10290,G10291,G10292,G10293,G10294,G10295,G10296,G10297,G10298,G10299,G10300,
       G10301,G10302,G10303,G10304,G10305,G10306,G10307,G10308,G10309,G10310,G10311,G10312,G10313,G10314,G10315,G10316,G10317,G10318,G10319,G10320,
       G10321,G10322,G10323,G10324,G10325,G10326,G10327,G10328,G10329,G10330,G10331,G10332,G10333,G10334,G10335,G10336,G10337,G10338,G10339,G10340,
       G10341,G10342,G10343,G10344,G10345,G10346,G10347,G10348,G10349,G10350,G10351,G10352,G10353,G10354,G10355,G10356,G10357,G10358,G10359,G10360,
       G10361,G10362,G10363,G10364,G10365,G10366,G10367,G10368,G10369,G10370,G10371,G10372,G10373,G10374,G10375,G10376,G10377,G10378,G10379,G10380,
       G10381,G10382,G10383,G10384,G10385,G10386,G10387,G10388,G10389,G10390,G10391,G10392,G10393,G10394,G10395,G10396,G10397,G10398,G10399,G10400,
       G10401,G10402,G10403,G10404,G10405,G10406,G10407,G10408,G10409,G10410,G10411,G10412,G10413,G10414,G10415,G10416,G10417,G10418,G10419,G10420,
       G10421,G10422,G10423,G10424,G10425,G10426,G10427,G10428,G10429,G10430,G10431,G10432,G10433,G10434,G10435,G10436,G10437,G10438,G10439,G10440,
       G10441,G10442,G10443,G10444,G10445,G10446,G10447,G10448,G10449,G10450,G10451,G10452,G10453,G10454,G10455,G10456,G10457,G10458,G10459,G10460,
       G10461,G10462,G10463,G10464,G10465,G10466,G10467,G10468,G10469,G10470,G10471,G10472,G10473,G10474,G10475,G10476,G10477,G10478,G10479,G10480,
       G10481,G10482,G10483,G10484,G10485,G10486,G10487,G10488,G10489,G10490,G10491,G10492,G10493,G10494,G10495,G10496,G10497,G10498,G10499,G10500,
       G10501,G10502,G10503,G10504,G10505,G10506,G10507,G10508,G10509,G10510,G10511,G10512,G10513,G10514,G10515,G10516,G10517,G10518,G10519,G10520,
       G10521,G10522,G10523,G10524,G10525,G10526,G10527,G10528,G10529,G10530,G10531,G10532,G10533,G10534,G10535,G10536,G10537,G10538,G10539,G10540,
       G10541,G10542,G10543,G10544,G10545,G10546,G10547,G10548,G10549,G10550,G10551,G10552,G10553,G10554,G10555,G10556,G10557,G10558,G10559,G10560,
       G10561,G10562,G10563,G10564,G10565,G10566,G10567,G10568,G10569,G10570,G10571,G10572,G10573,G10574,G10575,G10576,G10577,G10578,G10579,G10580,
       G10581,G10582,G10583,G10584,G10585,G10586,G10587,G10588,G10589,G10590,G10591,G10592,G10593,G10594,G10595,G10596,G10597,G10598,G10599,G10600,
       G10601,G10602,G10603,G10604,G10605,G10606,G10607,G10608,G10609,G10610,G10611,G10612,G10613,G10614,G10615,G10616,G10617,G10618,G10619,G10620,
       G10621,G10622,G10623,G10624,G10625,G10626,G10627,G10628,G10629,G10630,G10631,G10632,G10633,G10634,G10635,G10636,G10637,G10638,G10639,G10640,
       G10641,G10642,G10643,G10644,G10645,G10646,G10647,G10648,G10649,G10650,G10651,G10652,G10653,G10654,G10655,G10656,G10657,G10658,G10659,G10660,
       G10661,G10662,G10663,G10664,G10665,G10666,G10667,G10668,G10669,G10670,G10671,G10672,G10673,G10674,G10675,G10676,G10677,G10678,G10679,G10680,
       G10681,G10682,G10683,G10684,G10685,G10686,G10687,G10688,G10689,G10690,G10691,G10692,G10693,G10694,G10695,G10696,G10697,G10698,G10699,G10700,
       G10701,G10702,G10703,G10704,G10705,G10706,G10707,G10708,G10709,G10710,G10711,G10712,G10713,G10714,G10715,G10716,G10717,G10718,G10719,G10720,
       G10721,G10722,G10723,G10724,G10725,G10726,G10727,G10728,G10729,G10730,G10731,G10732,G10733,G10734,G10735,G10736,G10737,G10738,G10739,G10740,
       G10741,G10742,G10743,G10744,G10745,G10746,G10747,G10748,G10749,G10750,G10751,G10752,G10753,G10754,G10755,G10756,G10757,G10758,G10759,G10760,
       G10761,G10762,G10763,G10764,G10765,G10766,G10767,G10768,G10769,G10770,G10771,G10772,G10773,G10774,G10775,G10776,G10777,G10778,G10779,G10780,
       G10781,G10782,G10783,G10784,G10785,G10786,G10787,G10788,G10789,G10790,G10791,G10792,G10793,G10794,G10795,G10796,G10797,G10798,G10799,G10800,
       G10801,G10802,G10803,G10804,G10805,G10806,G10807,G10808,G10809,G10810,G10811,G10812,G10813,G10814,G10815,G10816,G10817,G10818,G10819,G10820,
       G10821,G10822,G10823,G10824,G10825,G10826,G10827,G10828,G10829,G10830,G10831,G10832,G10833,G10834,G10835,G10836,G10837,G10838,G10839,G10840,
       G10841,G10842,G10843,G10844,G10845,G10846,G10847,G10848,G10849,G10850,G10851,G10852,G10853,G10854,G10855,G10856,G10857,G10858,G10859,G10860,
       G10861,G10862,G10863,G10864,G10865,G10866,G10867,G10868,G10869,G10870,G10871,G10872,G10873,G10874,G10875,G10876,G10877,G10878,G10879,G10880,
       G10881,G10882,G10883,G10884,G10885,G10886,G10887,G10888,G10889,G10890,G10891,G10892,G10893,G10894,G10895,G10896,G10897,G10898,G10899,G10900,
       G10901,G10902,G10903,G10904,G10905,G10906,G10907,G10908,G10909,G10910,G10911,G10912,G10913,G10914,G10915,G10916,G10917,G10918,G10919,G10920,
       G10921,G10922,G10923,G10924,G10925,G10926,G10927,G10928,G10929,G10930,G10931,G10932,G10933,G10934,G10935,G10936,G10937,G10938,G10939,G10940,
       G10941,G10942,G10943,G10944,G10945,G10946,G10947,G10948,G10949,G10950,G10951,G10952,G10953,G10954,G10955,G10956,G10957,G10958,G10959,G10960,
       G10961,G10962,G10963,G10964,G10965,G10966,G10967,G10968,G10969,G10970,G10971,G10972,G10973,G10974,G10975,G10976,G10977,G10978,G10979,G10980,
       G10981,G10982,G10983,G10984,G10985,G10986,G10987,G10988,G10989,G10990,G10991,G10992,G10993,G10994,G10995,G10996,G10997,G10998,G10999,G11000,
       G11001,G11002,G11003,G11004,G11005,G11006,G11007,G11008,G11009,G11010,G11011,G11012,G11013,G11014,G11015,G11016,G11017,G11018,G11019,G11020,
       G11021,G11022,G11023,G11024,G11025,G11026,G11027,G11028,G11029,G11030,G11031,G11032,G11033,G11034,G11035,G11036,G11037,G11038,G11039,G11040,
       G11041,G11042,G11043,G11044,G11045,G11046,G11047,G11048,G11049,G11050,G11051,G11052,G11053,G11054,G11055,G11056,G11057,G11058,G11059,G11060,
       G11061,G11062,G11063,G11064,G11065,G11066,G11067,G11068,G11069,G11070,G11071,G11072,G11073,G11074,G11075,G11076,G11077,G11078,G11079,G11080,
       G11081,G11082,G11083,G11084,G11085,G11086,G11087,G11088,G11089,G11090,G11091,G11092,G11093,G11094,G11095,G11096,G11097,G11098,G11099,G11100,
       G11101,G11102,G11103,G11104,G11105,G11106,G11107,G11108,G11109,G11110,G11111,G11112,G11113,G11114,G11115,G11116,G11117,G11118,G11119,G11120,
       G11121,G11122,G11123,G11124,G11125,G11126,G11127,G11128,G11129,G11130,G11131,G11132,G11133,G11134,G11135,G11136,G11137,G11138,G11139,G11140,
       G11141,G11142,G11143,G11144,G11145,G11146,G11147,G11148,G11149,G11150,G11151,G11152,G11153,G11154,G11155,G11156,G11157,G11158,G11159,G11160,
       G11161,G11162,G11163,G11164,G11165,G11166,G11167,G11168,G11169,G11170,G11171,G11172,G11173,G11174,G11175,G11176,G11177,G11178,G11179,G11180,
       G11181,G11182,G11183,G11184,G11185,G11186,G11187,G11188,G11189,G11190,G11191,G11192,G11193,G11194,G11195,G11196,G11197,G11198,G11199,G11200,
       G11201,G11202,G11203,G11204,G11205,G11206,G11207,G11208,G11209,G11210,G11211,G11212,G11213,G11214,G11215,G11216,G11217,G11218,G11219,G11220,
       G11221,G11222,G11223,G11224,G11225,G11226,G11227,G11228,G11229,G11230,G11231,G11232,G11233,G11234,G11235,G11236,G11237,G11238,G11239,G11240,
       G11241,G11242,G11243,G11244,G11245,G11246,G11247,G11248,G11249,G11250,G11251,G11252,G11253,G11254,G11255,G11256,G11257,G11258,G11259,G11260,
       G11261,G11262,G11263,G11264,G11265,G11266,G11267,G11268,G11269,G11270,G11271,G11272,G11273,G11274,G11275,G11276,G11277,G11278,G11279,G11280,
       G11281,G11282,G11283,G11284,G11285,G11286,G11287,G11288,G11289,G11290,G11291,G11292,G11293,G11294,G11295,G11296,G11297,G11298,G11299,G11300,
       G11301,G11302,G11303,G11304,G11305,G11306,G11307,G11308,G11309,G11310,G11311,G11312,G11313,G11314,G11315,G11316,G11317,G11318,G11319,G11320,
       G11321,G11322,G11323,G11324,G11325,G11326,G11327,G11328,G11329,G11330,G11331,G11332,G11333,G11334,G11335,G11336,G11337,G11338,G11339,G11340,
       G11341,G11342,G11343,G11344,G11345,G11346,G11347,G11348,G11349,G11350,G11351,G11352,G11353,G11354,G11355,G11356,G11357,G11358,G11359,G11360,
       G11361,G11362,G11363,G11364,G11365,G11366,G11367,G11368,G11369,G11370,G11371,G11372,G11373,G11374,G11375,G11376,G11377,G11378,G11379,G11380,
       G11381,G11382,G11383,G11384,G11385,G11386,G11387,G11388,G11389,G11390,G11391,G11392,G11393,G11394,G11395,G11396,G11397,G11398,G11399,G11400,
       G11401,G11402,G11403,G11404,G11405,G11406,G11407,G11408,G11409,G11410,G11411,G11412,G11413,G11414,G11415,G11416,G11417,G11418,G11419,G11420,
       G11421,G11422,G11423,G11424,G11425,G11426,G11427,G11428,G11429,G11430,G11431,G11432,G11433,G11434,G11435,G11436,G11437,G11438,G11439,G11440,
       G11441,G11442,G11443,G11444,G11445,G11446,G11447,G11448,G11449,G11450,G11451,G11452,G11453,G11454,G11455,G11456,G11457,G11458,G11459,G11460,
       G11461,G11462,G11463,G11464,G11465,G11466,G11467,G11468,G11469,G11470,G11471,G11472,G11473,G11474,G11475,G11476,G11477,G11478,G11479,G11480,
       G11481,G11482,G11483,G11484,G11485,G11486,G11487,G11488,G11489,G11490,G11491,G11492,G11493,G11494,G11495,G11496,G11497,G11498,G11499,G11500,
       G11501,G11502,G11503,G11504,G11505,G11506,G11507,G11508,G11509,G11510,G11511,G11512,G11513,G11514,G11515,G11516,G11517,G11518,G11519,G11520,
       G11521,G11522,G11523,G11524,G11525,G11526,G11527,G11528,G11529,G11530,G11531,G11532,G11533,G11534,G11535,G11536,G11537,G11538,G11539,G11540,
       G11541,G11542,G11543,G11544,G11545,G11546,G11547,G11548,G11549,G11550,G11551,G11552,G11553,G11554,G11555,G11556,G11557,G11558,G11559,G11560,
       G11561,G11562,G11563,G11564,G11565,G11566,G11567,G11568,G11569,G11570,G11571,G11572,G11573,G11574,G11575,G11576,G11577,G11578,G11579,G11580,
       G11581,G11582,G11583,G11584,G11585,G11586,G11587,G11588,G11589,G11590,G11591,G11592,G11593,G11594,G11595,G11596,G11597,G11598,G11599,G11600,
       G11601,G11602,G11603,G11604,G11605,G11606,G11607,G11608,G11609,G11610,G11611,G11612,G11613,G11614,G11615,G11616,G11617,G11618,G11619,G11620,
       G11621,G11622,G11623,G11624,G11625,G11626,G11627,G11628,G11629,G11630,G11631,G11632,G11633,G11634,G11635,G11636,G11637,G11638,G11639,G11640,
       G11641,G11642,G11643,G11644,G11645,G11646,G11647,G11648,G11649,G11650,G11651,G11652,G11653,G11654,G11655,G11656,G11657,G11658,G11659,G11660,
       G11661,G11662,G11663,G11664,G11665,G11666,G11667,G11668,G11669,G11670,G11671,G11672,G11673,G11674,G11675,G11676,G11677,G11678,G11679,G11680,
       G11681,G11682,G11683,G11684,G11685,G11686,G11687,G11688,G11689,G11690,G11691,G11692,G11693,G11694,G11695,G11696,G11697,G11698,G11699,G11700,
       G11701,G11702,G11703,G11704,G11705,G11706,G11707,G11708,G11709,G11710,G11711,G11712,G11713,G11714,G11715,G11716,G11717,G11718,G11719,G11720,
       G11721,G11722,G11723,G11724,G11725,G11726,G11727,G11728,G11729,G11730,G11731,G11732,G11733,G11734,G11735,G11736,G11737,G11738,G11739,G11740,
       G11741,G11742,G11743,G11744,G11745,G11746,G11747,G11748,G11749,G11750,G11751,G11752,G11753,G11754,G11755,G11756,G11757,G11758,G11759,G11760,
       G11761,G11762,G11763,G11764,G11765,G11766,G11767,G11768,G11769,G11770,G11771,G11772,G11773,G11774,G11775,G11776,G11777,G11778,G11779,G11780,
       G11781,G11782,G11783,G11784,G11785,G11786,G11787,G11788,G11789,G11790,G11791,G11792,G11793,G11794,G11795,G11796,G11797,G11798,G11799,G11800,
       G11801,G11802,G11803,G11804,G11805,G11806,G11807,G11808,G11809,G11810,G11811,G11812,G11813,G11814,G11815,G11816,G11817,G11818,G11819,G11820,
       G11821,G11822,G11823,G11824,G11825,G11826,G11827,G11828,G11829,G11830,G11831,G11832,G11833,G11834,G11835,G11836,G11837,G11838,G11839,G11840,
       G11841,G11842,G11843,G11844,G11845,G11846,G11847,G11848,G11849,G11850,G11851,G11852,G11853,G11854,G11855,G11856,G11857,G11858,G11859,G11860,
       G11861,G11862,G11863,G11864,G11865,G11866,G11867,G11868,G11869,G11870,G11871,G11872,G11873,G11874,G11875,G11876,G11877,G11878,G11879,G11880,
       G11881,G11882,G11883,G11884,G11885,G11886,G11887,G11888,G11889,G11890,G11891,G11892,G11893,G11894,G11895,G11896,G11897,G11898,G11899,G11900,
       G11901,G11902,G11903,G11904,G11905,G11906,G11907,G11908,G11909,G11910,G11911,G11912,G11913,G11914,G11915,G11916,G11917,G11918,G11919,G11920,
       G11921,G11922,G11923,G11924,G11925,G11926,G11927,G11928,G11929,G11930,G11931,G11932,G11933,G11934,G11935,G11936,G11937,G11938,G11939,G11940,
       G11941,G11942,G11943,G11944,G11945,G11946,G11947,G11948,G11949,G11950,G11951,G11952,G11953,G11954,G11955,G11956,G11957,G11958,G11959,G11960,
       G11961,G11962,G11963,G11964,G11965,G11966,G11967,G11968,G11969,G11970,G11971,G11972,G11973,G11974,G11975,G11976,G11977,G11978,G11979,G11980,
       G11981,G11982,G11983,G11984,G11985,G11986,G11987,G11988,G11989,G11990,G11991,G11992,G11993,G11994,G11995,G11996,G11997,G11998,G11999,G12000,
       G12001,G12002,G12003,G12004,G12005,G12006,G12007,G12008,G12009,G12010,G12011,G12012,G12013,G12014,G12015,G12016,G12017,G12018,G12019,G12020,
       G12021,G12022,G12023,G12024,G12025,G12026,G12027,G12028,G12029,G12030,G12031,G12032,G12033,G12034,G12035,G12036,G12037,G12038,G12039,G12040,
       G12041,G12042,G12043,G12044,G12045,G12046,G12047,G12048,G12049,G12050,G12051,G12052,G12053,G12054,G12055,G12056,G12057,G12058,G12059,G12060,
       G12061,G12062,G12063,G12064,G12065,G12066,G12067,G12068,G12069,G12070,G12071,G12072,G12073,G12074,G12075,G12076,G12077,G12078,G12079,G12080,
       G12081,G12082,G12083,G12084,G12085,G12086,G12087,G12088,G12089,G12090,G12091,G12092,G12093,G12094,G12095,G12096,G12097,G12098,G12099,G12100,
       G12101,G12102,G12103,G12104,G12105,G12106,G12107,G12108,G12109,G12110,G12111,G12112,G12113,G12114,G12115,G12116,G12117,G12118,G12119,G12120,
       G12121,G12122,G12123,G12124,G12125,G12126,G12127,G12128,G12129,G12130,G12131,G12132,G12133,G12134,G12135,G12136,G12137,G12138,G12139,G12140,
       G12141,G12142,G12143,G12144,G12145,G12146,G12147,G12148,G12149,G12150,G12151,G12152,G12153,G12154,G12155,G12156,G12157,G12158,G12159,G12160,
       G12161,G12162,G12163,G12164,G12165,G12166,G12167,G12168,G12169,G12170,G12171,G12172,G12173,G12174,G12175,G12176,G12177,G12178,G12179,G12180,
       G12181,G12182,G12183,G12184,G12185,G12186,G12187,G12188,G12189,G12190,G12191,G12192,G12193,G12194,G12195,G12196,G12197,G12198,G12199,G12200,
       G12201,G12202,G12203,G12204,G12205,G12206,G12207,G12208,G12209,G12210,G12211,G12212,G12213,G12214,G12215,G12216,G12217,G12218,G12219,G12220,
       G12221,G12222,G12223,G12224,G12225,G12226,G12227,G12228,G12229,G12230,G12231,G12232,G12233,G12234,G12235,G12236,G12237,G12238,G12239,G12240,
       G12241,G12242,G12243,G12244,G12245,G12246,G12247,G12248,G12249,G12250,G12251,G12252,G12253,G12254,G12255,G12256,G12257,G12258,G12259,G12260,
       G12261,G12262,G12263,G12264,G12265,G12266,G12267,G12268,G12269,G12270,G12271,G12272,G12273,G12274,G12275,G12276,G12277,G12278,G12279,G12280,
       G12281,G12282,G12283,G12284,G12285,G12286,G12287,G12288,G12289,G12290,G12291,G12292,G12293,G12294,G12295,G12296,G12297,G12298,G12299,G12300,
       G12301,G12302,G12303,G12304,G12305,G12306,G12307,G12308,G12309,G12310,G12311,G12312,G12313,G12314,G12315,G12316,G12317,G12318,G12319,G12320,
       G12321,G12322,G12323,G12324,G12325,G12326,G12327,G12328,G12329,G12330,G12331,G12332,G12333,G12334,G12335,G12336,G12337,G12338,G12339,G12340,
       G12341,G12342,G12343,G12344,G12345,G12346,G12347,G12348,G12349,G12350,G12351,G12352,G12353,G12354,G12355,G12356,G12357,G12358,G12359,G12360,
       G12361,G12362,G12363,G12364,G12365,G12366,G12367,G12368,G12369,G12370,G12371,G12372,G12373,G12374,G12375,G12376,G12377,G12378,G12379,G12380,
       G12381,G12382,G12383,G12384,G12385,G12386,G12387,G12388,G12389,G12390,G12391,G12392,G12393,G12394,G12395,G12396,G12397,G12398,G12399,G12400,
       G12401,G12402,G12403,G12404,G12405,G12406,G12407,G12408,G12409,G12410,G12411,G12412,G12413,G12414,G12415,G12416,G12417,G12418,G12419,G12420,
       G12421,G12422,G12423,G12424,G12425,G12426,G12427,G12428,G12429,G12430,G12431,G12432,G12433,G12434,G12435,G12436,G12437,G12438,G12439,G12440,
       G12441,G12442,G12443,G12444,G12445,G12446,G12447,G12448,G12449,G12450,G12451,G12452,G12453,G12454,G12455,G12456,G12457,G12458,G12459,G12460,
       G12461,G12462,G12463,G12464,G12465,G12466,G12467,G12468,G12469,G12470,G12471,G12472,G12473,G12474,G12475,G12476,G12477,G12478,G12479,G12480,
       G12481,G12482,G12483,G12484,G12485,G12486,G12487,G12488,G12489,G12490,G12491,G12492,G12493,G12494,G12495,G12496,G12497,G12498,G12499,G12500,
       G12501,G12502,G12503,G12504,G12505,G12506,G12507,G12508,G12509,G12510,G12511,G12512,G12513,G12514,G12515,G12516,G12517,G12518,G12519,G12520,
       G12521,G12522,G12523,G12524,G12525,G12526,G12527,G12528,G12529,G12530,G12531,G12532,G12533,G12534,G12535,G12536,G12537,G12538,G12539,G12540,
       G12541,G12542,G12543,G12544,G12545,G12546,G12547,G12548,G12549,G12550,G12551,G12552,G12553,G12554,G12555,G12556,G12557,G12558,G12559,G12560,
       G12561,G12562,G12563,G12564,G12565,G12566,G12567,G12568,G12569,G12570,G12571,G12572,G12573,G12574,G12575,G12576,G12577,G12578,G12579,G12580,
       G12581,G12582,G12583,G12584,G12585,G12586,G12587,G12588,G12589,G12590,G12591,G12592,G12593,G12594,G12595,G12596,G12597,G12598,G12599,G12600,
       G12601,G12602,G12603,G12604,G12605,G12606,G12607,G12608,G12609,G12610,G12611,G12612,G12613,G12614,G12615,G12616,G12617,G12618,G12619,G12620,
       G12621,G12622,G12623,G12624,G12625,G12626,G12627,G12628,G12629,G12630,G12631,G12632,G12633,G12634,G12635,G12636,G12637,G12638,G12639,G12640,
       G12641,G12642,G12643,G12644,G12645,G12646,G12647,G12648,G12649,G12650,G12651,G12652,G12653,G12654,G12655,G12656,G12657,G12658,G12659,G12660,
       G12661,G12662,G12663,G12664,G12665,G12666,G12667,G12668,G12669,G12670,G12671,G12672,G12673,G12674,G12675,G12676,G12677,G12678,G12679,G12680,
       G12681,G12682,G12683,G12684,G12685,G12686,G12687,G12688,G12689,G12690,G12691,G12692,G12693,G12694,G12695,G12696,G12697,G12698,G12699,G12700,
       G12701,G12702,G12703,G12704,G12705,G12706,G12707,G12708,G12709,G12710,G12711,G12712,G12713,G12714,G12715,G12716,G12717,G12718,G12719,G12720,
       G12721,G12722,G12723,G12724,G12725,G12726,G12727,G12728,G12729,G12730,G12731,G12732,G12733,G12734,G12735,G12736,G12737,G12738,G12739,G12740,
       G12741,G12742,G12743,G12744,G12745,G12746,G12747,G12748,G12749,G12750,G12751,G12752,G12753,G12754,G12755,G12756,G12757,G12758,G12759,G12760,
       G12761,G12762,G12763,G12764,G12765,G12766,G12767,G12768,G12769,G12770,G12771,G12772,G12773,G12774,G12775,G12776,G12777,G12778,G12779,G12780,
       G12781,G12782,G12783,G12784,G12785,G12786,G12787,G12788,G12789,G12790,G12791,G12792,G12793,G12794,G12795,G12796,G12797,G12798,G12799,G12800,
       G12801,G12802,G12803,G12804,G12805,G12806,G12807,G12808,G12809,G12810,G12811,G12812,G12813,G12814,G12815,G12816,G12817,G12818,G12819,G12820,
       G12821,G12822,G12823,G12824,G12825,G12826,G12827,G12828,G12829,G12830,G12831,G12832,G12833,G12834,G12835,G12836,G12837,G12838,G12839,G12840,
       G12841,G12842,G12843,G12844,G12845,G12846,G12847,G12848,G12849,G12850,G12851,G12852,G12853,G12854,G12855,G12856,G12857,G12858,G12859,G12860,
       G12861,G12862,G12863,G12864,G12865,G12866,G12867,G12868,G12869,G12870,G12871,G12872,G12873,G12874,G12875,G12876,G12877,G12878,G12879,G12880,
       G12881,G12882,G12883,G12884,G12885,G12886,G12887,G12888,G12889,G12890,G12891,G12892,G12893,G12894,G12895,G12896,G12897,G12898,G12899,G12900,
       G12901,G12902,G12903,G12904,G12905,G12906,G12907,G12908,G12909,G12910,G12911,G12912,G12913,G12914,G12915,G12916,G12917,G12918,G12919,G12920,
       G12921,G12922,G12923,G12924,G12925,G12926,G12927,G12928,G12929,G12930,G12931,G12932,G12933,G12934,G12935,G12936,G12937,G12938,G12939,G12940,
       G12941,G12942,G12943,G12944,G12945,G12946,G12947,G12948,G12949,G12950,G12951,G12952,G12953,G12954,G12955,G12956,G12957,G12958,G12959,G12960,
       G12961,G12962,G12963,G12964,G12965,G12966,G12967,G12968,G12969,G12970,G12971,G12972,G12973,G12974,G12975,G12976,G12977,G12978,G12979,G12980,
       G12981,G12982,G12983,G12984,G12985,G12986,G12987,G12988,G12989,G12990,G12991,G12992,G12993,G12994,G12995,G12996,G12997,G12998,G12999,G13000,
       G13001,G13002,G13003,G13004,G13005,G13006,G13007,G13008,G13009,G13010,G13011,G13012,G13013,G13014,G13015,G13016,G13017,G13018,G13019,G13020,
       G13021,G13022,G13023,G13024,G13025,G13026,G13027,G13028,G13029,G13030,G13031,G13032,G13033,G13034,G13035,G13036,G13037,G13038,G13039,G13040,
       G13041,G13042,G13043,G13044,G13045,G13046,G13047,G13048,G13049,G13050,G13051,G13052,G13053,G13054,G13055,G13056,G13057,G13058,G13059,G13060,
       G13061,G13062,G13063,G13064,G13065,G13066,G13067,G13068,G13069,G13070,G13071,G13072,G13073,G13074,G13075,G13076,G13077,G13078,G13079,G13080,
       G13081,G13082,G13083,G13084,G13085,G13086,G13087,G13088,G13089,G13090,G13091,G13092,G13093,G13094,G13095,G13096,G13097,G13098,G13099,G13100,
       G13101,G13102,G13103,G13104,G13105,G13106,G13107,G13108,G13109,G13110,G13111,G13112,G13113,G13114,G13115,G13116,G13117,G13118,G13119,G13120,
       G13121,G13122,G13123,G13124,G13125,G13126,G13127,G13128,G13129,G13130,G13131,G13132,G13133,G13134,G13135,G13136,G13137,G13138,G13139,G13140,
       G13141,G13142,G13143,G13144,G13145,G13146,G13147,G13148,G13149,G13150,G13151,G13152,G13153,G13154,G13155,G13156,G13157,G13158,G13159,G13160,
       G13161,G13162,G13163,G13164,G13165,G13166,G13167,G13168,G13169,G13170,G13171,G13172,G13173,G13174,G13175,G13176,G13177,G13178,G13179,G13180,
       G13181,G13182,G13183,G13184,G13185,G13186,G13187,G13188,G13189,G13190,G13191,G13192,G13193,G13194,G13195,G13196,G13197,G13198,G13199,G13200,
       G13201,G13202,G13203,G13204,G13205,G13206,G13207,G13208,G13209,G13210,G13211,G13212,G13213,G13214,G13215,G13216,G13217,G13218,G13219,G13220,
       G13221,G13222,G13223,G13224,G13225,G13226,G13227,G13228,G13229,G13230,G13231,G13232,G13233,G13234,G13235,G13236,G13237,G13238,G13239,G13240,
       G13241,G13242,G13243,G13244,G13245,G13246,G13247,G13248,G13249,G13250,G13251,G13252,G13253,G13254,G13255,G13256,G13257,G13258,G13259,G13260,
       G13261,G13262,G13263,G13264,G13265,G13266,G13267,G13268,G13269,G13270,G13271,G13272,G13273,G13274,G13275,G13276,G13277,G13278,G13279,G13280,
       G13281,G13282,G13283,G13284,G13285,G13286,G13287,G13288,G13289,G13290,G13291,G13292,G13293,G13294,G13295,G13296,G13297,G13298,G13299,G13300,
       G13301,G13302,G13303,G13304,G13305,G13306,G13307,G13308,G13309,G13310,G13311,G13312,G13313,G13314,G13315,G13316,G13317,G13318,G13319,G13320,
       G13321,G13322,G13323,G13324,G13325,G13326,G13327,G13328,G13329,G13330,G13331,G13332,G13333,G13334,G13335,G13336,G13337,G13338,G13339,G13340,
       G13341,G13342,G13343,G13344,G13345,G13346,G13347,G13348,G13349,G13350,G13351,G13352,G13353,G13354,G13355,G13356,G13357,G13358,G13359,G13360,
       G13361,G13362,G13363,G13364,G13365,G13366,G13367,G13368,G13369,G13370,G13371,G13372,G13373,G13374,G13375,G13376,G13377,G13378,G13379,G13380,
       G13381,G13382,G13383,G13384,G13385,G13386,G13387,G13388,G13389,G13390,G13391,G13392,G13393,G13394,G13395,G13396,G13397,G13398,G13399,G13400,
       G13401,G13402,G13403,G13404,G13405,G13406,G13407,G13408,G13409,G13410,G13411,G13412,G13413,G13414,G13415,G13416,G13417,G13418,G13419,G13420,
       G13421,G13422,G13423,G13424,G13425,G13426,G13427,G13428,G13429,G13430,G13431,G13432,G13433,G13434,G13435,G13436,G13437,G13438,G13439,G13440,
       G13441,G13442,G13443,G13444,G13445,G13446,G13447,G13448,G13449,G13450,G13451,G13452,G13453,G13454,G13455,G13456,G13457,G13458,G13459,G13460,
       G13461,G13462,G13463,G13464,G13465,G13466,G13467,G13468,G13469,G13470,G13471,G13472,G13473,G13474,G13475,G13476,G13477,G13478,G13479,G13480,
       G13481,G13482,G13483,G13484,G13485,G13486,G13487,G13488,G13489,G13490,G13491,G13492,G13493,G13494,G13495,G13496,G13497,G13498,G13499,G13500,
       G13501,G13502,G13503,G13504,G13505,G13506,G13507,G13508,G13509,G13510,G13511,G13512,G13513,G13514,G13515,G13516,G13517,G13518,G13519,G13520,
       G13521,G13522,G13523,G13524,G13525,G13526,G13527,G13528,G13529,G13530,G13531,G13532,G13533,G13534,G13535,G13536,G13537,G13538,G13539,G13540,
       G13541,G13542,G13543,G13544,G13545,G13546,G13547,G13548,G13549,G13550,G13551,G13552,G13553,G13554,G13555,G13556,G13557,G13558,G13559,G13560,
       G13561,G13562,G13563,G13564,G13565,G13566,G13567,G13568,G13569,G13570,G13571,G13572,G13573,G13574,G13575,G13576,G13577,G13578,G13579,G13580,
       G13581,G13582,G13583,G13584,G13585,G13586,G13587,G13588,G13589,G13590,G13591,G13592,G13593,G13594,G13595,G13596,G13597,G13598,G13599,G13600,
       G13601,G13602,G13603,G13604,G13605,G13606,G13607,G13608,G13609,G13610,G13611,G13612,G13613,G13614,G13615,G13616,G13617,G13618,G13619,G13620,
       G13621,G13622,G13623,G13624,G13625,G13626,G13627,G13628,G13629,G13630,G13631,G13632,G13633,G13634,G13635,G13636,G13637,G13638,G13639,G13640,
       G13641,G13642,G13643,G13644,G13645,G13646,G13647,G13648,G13649,G13650,G13651,G13652,G13653,G13654,G13655,G13656,G13657,G13658,G13659,G13660,
       G13661,G13662,G13663,G13664,G13665,G13666,G13667,G13668,G13669,G13670,G13671,G13672,G13673,G13674,G13675,G13676,G13677,G13678,G13679,G13680,
       G13681,G13682,G13683,G13684,G13685,G13686,G13687,G13688,G13689,G13690,G13691,G13692,G13693,G13694,G13695,G13696,G13697,G13698,G13699,G13700,
       G13701,G13702,G13703,G13704,G13705,G13706,G13707,G13708,G13709,G13710,G13711,G13712,G13713,G13714,G13715,G13716,G13717,G13718,G13719,G13720,
       G13721,G13722,G13723,G13724,G13725,G13726,G13727,G13728,G13729,G13730,G13731,G13732,G13733,G13734,G13735,G13736,G13737,G13738,G13739,G13740,
       G13741,G13742,G13743,G13744,G13745,G13746,G13747,G13748,G13749,G13750,G13751,G13752,G13753,G13754,G13755,G13756,G13757,G13758,G13759,G13760,
       G13761,G13762,G13763,G13764,G13765,G13766,G13767,G13768,G13769,G13770,G13771,G13772,G13773,G13774,G13775,G13776,G13777,G13778,G13779,G13780,
       G13781,G13782,G13783,G13784,G13785,G13786,G13787,G13788,G13789,G13790,G13791,G13792,G13793,G13794,G13795,G13796,G13797,G13798,G13799,G13800,
       G13801,G13802,G13803,G13804,G13805,G13806,G13807,G13808,G13809,G13810,G13811,G13812,G13813,G13814,G13815,G13816,G13817,G13818,G13819,G13820,
       G13821,G13822,G13823,G13824,G13825,G13826,G13827,G13828,G13829,G13830,G13831,G13832,G13833,G13834,G13835,G13836,G13837,G13838,G13839,G13840,
       G13841,G13842,G13843,G13844,G13845,G13846,G13847,G13848,G13849,G13850,G13851,G13852,G13853,G13854,G13855,G13856,G13857,G13858,G13859,G13860,
       G13861,G13862,G13863,G13864,G13865,G13866,G13867,G13868,G13869,G13870,G13871,G13872,G13873,G13874,G13875,G13876,G13877,G13878,G13879,G13880,
       G13881,G13882,G13883,G13884,G13885,G13886,G13887,G13888,G13889,G13890,G13891,G13892,G13893,G13894,G13895,G13896,G13897,G13898,G13899,G13900,
       G13901,G13902,G13903,G13904,G13905,G13906,G13907,G13908,G13909,G13910,G13911,G13912,G13913,G13914,G13915,G13916,G13917,G13918,G13919,G13920,
       G13921,G13922,G13923,G13924,G13925,G13926,G13927,G13928,G13929,G13930,G13931,G13932,G13933,G13934,G13935,G13936,G13937,G13938,G13939,G13940,
       G13941,G13942,G13943,G13944,G13945,G13946,G13947,G13948,G13949,G13950,G13951,G13952,G13953,G13954,G13955,G13956,G13957,G13958,G13959,G13960,
       G13961,G13962,G13963,G13964,G13965,G13966,G13967,G13968,G13969,G13970,G13971,G13972,G13973,G13974,G13975,G13976,G13977,G13978,G13979,G13980,
       G13981,G13982,G13983,G13984,G13985,G13986,G13987,G13988,G13989,G13990,G13991,G13992,G13993,G13994,G13995,G13996,G13997,G13998,G13999,G14000,
       G14001,G14002,G14003,G14004,G14005,G14006,G14007,G14008,G14009,G14010,G14011,G14012,G14013,G14014,G14015,G14016,G14017,G14018,G14019,G14020,
       G14021,G14022,G14023,G14024,G14025,G14026,G14027,G14028,G14029,G14030,G14031,G14032,G14033,G14034,G14035,G14036,G14037,G14038,G14039,G14040,
       G14041,G14042,G14043,G14044,G14045,G14046,G14047,G14048,G14049,G14050,G14051,G14052,G14053,G14054,G14055,G14056,G14057,G14058,G14059,G14060,
       G14061,G14062,G14063,G14064,G14065,G14066,G14067,G14068,G14069,G14070,G14071,G14072,G14073,G14074,G14075,G14076,G14077,G14078,G14079,G14080,
       G14081,G14082,G14083,G14084,G14085,G14086,G14087,G14088,G14089,G14090,G14091,G14092,G14093,G14094,G14095,G14096,G14097,G14098,G14099,G14100,
       G14101,G14102,G14103,G14104,G14105,G14106,G14107,G14108,G14109,G14110,G14111,G14112,G14113,G14114,G14115,G14116,G14117,G14118,G14119,G14120,
       G14121,G14122,G14123,G14124,G14125,G14126,G14127,G14128,G14129,G14130,G14131,G14132,G14133,G14134,G14135,G14136,G14137,G14138,G14139,G14140,
       G14141,G14142,G14143,G14144,G14145,G14146,G14147,G14148,G14149,G14150,G14151,G14152,G14153,G14154,G14155,G14156,G14157,G14158,G14159,G14160,
       G14161,G14162,G14163,G14164,G14165,G14166,G14167,G14168,G14169,G14170,G14171,G14172,G14173,G14174,G14175,G14176,G14177,G14178,G14179,G14180,
       G14181,G14182,G14183,G14184,G14185,G14186,G14187,G14188,G14189,G14190,G14191,G14192,G14193,G14194,G14195,G14196,G14197,G14198,G14199,G14200,
       G14201,G14202,G14203,G14204,G14205,G14206,G14207,G14208,G14209,G14210,G14211,G14212,G14213,G14214,G14215,G14216,G14217,G14218,G14219,G14220,
       G14221,G14222,G14223,G14224,G14225,G14226,G14227,G14228,G14229,G14230,G14231,G14232,G14233,G14234,G14235,G14236,G14237,G14238,G14239,G14240,
       G14241,G14242,G14243,G14244,G14245,G14246,G14247,G14248,G14249,G14250,G14251,G14252,G14253,G14254,G14255,G14256,G14257,G14258,G14259,G14260,
       G14261,G14262,G14263,G14264,G14265,G14266,G14267,G14268,G14269,G14270,G14271,G14272,G14273,G14274,G14275,G14276,G14277,G14278,G14279,G14280,
       G14281,G14282,G14283,G14284,G14285,G14286,G14287,G14288,G14289,G14290,G14291,G14292,G14293,G14294,G14295,G14296,G14297,G14298,G14299,G14300,
       G14301,G14302,G14303,G14304,G14305,G14306,G14307,G14308,G14309,G14310,G14311,G14312,G14313,G14314,G14315,G14316,G14317,G14318,G14319,G14320,
       G14321,G14322,G14323,G14324,G14325,G14326,G14327,G14328,G14329,G14330,G14331,G14332,G14333,G14334,G14335,G14336,G14337,G14338,G14339,G14340,
       G14341,G14342,G14343,G14344,G14345,G14346,G14347,G14348,G14349,G14350,G14351,G14352,G14353,G14354,G14355,G14356,G14357,G14358,G14359,G14360,
       G14361,G14362,G14363,G14364,G14365,G14366,G14367,G14368,G14369,G14370,G14371,G14372,G14373,G14374,G14375,G14376,G14377,G14378,G14379,G14380,
       G14381,G14382,G14383,G14384,G14385,G14386,G14387,G14388,G14389,G14390,G14391,G14392,G14393,G14394,G14395,G14396,G14397,G14398,G14399,G14400,
       G14401,G14402,G14403,G14404,G14405,G14406,G14407,G14408,G14409,G14410,G14411,G14412,G14413,G14414,G14415,G14416,G14417,G14418,G14419,G14420,
       G14421,G14422,G14423,G14424,G14425,G14426,G14427,G14428,G14429,G14430,G14431,G14432,G14433,G14434,G14435,G14436,G14437,G14438,G14439,G14440,
       G14441,G14442,G14443,G14444,G14445,G14446,G14447,G14448,G14449,G14450,G14451,G14452,G14453,G14454,G14455,G14456,G14457,G14458,G14459,G14460,
       G14461,G14462,G14463,G14464,G14465,G14466,G14467,G14468,G14469,G14470,G14471,G14472,G14473,G14474,G14475,G14476,G14477,G14478,G14479,G14480,
       G14481,G14482,G14483,G14484,G14485,G14486,G14487,G14488,G14489,G14490,G14491,G14492,G14493,G14494,G14495,G14496,G14497,G14498,G14499,G14500,
       G14501,G14502,G14503,G14504,G14505,G14506,G14507,G14508,G14509,G14510,G14511,G14512,G14513,G14514,G14515,G14516,G14517,G14518,G14519,G14520,
       G14521,G14522,G14523,G14524,G14525,G14526,G14527,G14528,G14529,G14530,G14531,G14532,G14533,G14534,G14535,G14536,G14537,G14538,G14539,G14540,
       G14541,G14542,G14543,G14544,G14545,G14546,G14547,G14548,G14549,G14550,G14551,G14552,G14553,G14554,G14555,G14556,G14557,G14558,G14559,G14560,
       G14561,G14562,G14563,G14564,G14565,G14566,G14567,G14568,G14569,G14570,G14571,G14572,G14573,G14574,G14575,G14576,G14577,G14578,G14579,G14580,
       G14581,G14582,G14583,G14584,G14585,G14586,G14587,G14588,G14589,G14590,G14591,G14592,G14593,G14594,G14595,G14596,G14597,G14598,G14599,G14600,
       G14601,G14602,G14603,G14604,G14605,G14606,G14607,G14608,G14609,G14610,G14611,G14612,G14613,G14614,G14615,G14616,G14617,G14618,G14619,G14620,
       G14621,G14622,G14623,G14624,G14625,G14626,G14627,G14628,G14629,G14630,G14631,G14632,G14633,G14634,G14635,G14636,G14637,G14638,G14639,G14640,
       G14641,G14642,G14643,G14644,G14645,G14646,G14647,G14648,G14649,G14650,G14651,G14652,G14653,G14654,G14655,G14656,G14657,G14658,G14659,G14660,
       G14661,G14662,G14663,G14664,G14665,G14666,G14667,G14668,G14669,G14670,G14671,G14672,G14673,G14674,G14675,G14676,G14677,G14678,G14679,G14680,
       G14681,G14682,G14683,G14684,G14685,G14686,G14687,G14688,G14689,G14690,G14691,G14692,G14693,G14694,G14695,G14696,G14697,G14698,G14699,G14700,
       G14701,G14702,G14703,G14704,G14705,G14706,G14707,G14708,G14709,G14710,G14711,G14712,G14713,G14714,G14715,G14716,G14717,G14718,G14719,G14720,
       G14721,G14722,G14723,G14724,G14725,G14726,G14727,G14728,G14729,G14730,G14731,G14732,G14733,G14734,G14735,G14736,G14737,G14738,G14739,G14740,
       G14741,G14742,G14743,G14744,G14745,G14746,G14747,G14748,G14749,G14750,G14751,G14752,G14753,G14754,G14755,G14756,G14757,G14758,G14759,G14760,
       G14761,G14762,G14763,G14764,G14765,G14766,G14767,G14768,G14769,G14770,G14771,G14772,G14773,G14774,G14775,G14776,G14777,G14778,G14779,G14780,
       G14781,G14782,G14783,G14784,G14785,G14786,G14787,G14788,G14789,G14790,G14791,G14792,G14793,G14794,G14795,G14796,G14797,G14798,G14799,G14800,
       G14801,G14802,G14803,G14804,G14805,G14806,G14807,G14808,G14809,G14810,G14811,G14812,G14813,G14814,G14815,G14816,G14817,G14818,G14819,G14820,
       G14821,G14822,G14823,G14824,G14825,G14826,G14827,G14828,G14829,G14830,G14831,G14832,G14833,G14834,G14835,G14836,G14837,G14838,G14839,G14840,
       G14841,G14842,G14843,G14844,G14845,G14846,G14847,G14848,G14849,G14850,G14851,G14852,G14853,G14854,G14855,G14856,G14857,G14858,G14859,G14860,
       G14861,G14862,G14863,G14864,G14865,G14866,G14867,G14868,G14869,G14870,G14871,G14872,G14873,G14874,G14875,G14876,G14877,G14878,G14879,G14880,
       G14881,G14882,G14883,G14884,G14885,G14886,G14887,G14888,G14889,G14890,G14891,G14892,G14893,G14894,G14895,G14896,G14897,G14898,G14899,G14900,
       G14901,G14902,G14903,G14904,G14905,G14906,G14907,G14908,G14909,G14910,G14911,G14912,G14913,G14914,G14915,G14916,G14917,G14918,G14919,G14920,
       G14921,G14922,G14923,G14924,G14925,G14926,G14927,G14928,G14929,G14930,G14931,G14932,G14933,G14934,G14935,G14936,G14937,G14938,G14939,G14940,
       G14941,G14942,G14943,G14944,G14945,G14946,G14947,G14948,G14949,G14950,G14951,G14952,G14953,G14954,G14955,G14956,G14957,G14958,G14959,G14960,
       G14961,G14962,G14963,G14964,G14965,G14966,G14967,G14968,G14969,G14970,G14971,G14972,G14973,G14974,G14975,G14976,G14977,G14978,G14979,G14980,
       G14981,G14982,G14983,G14984,G14985,G14986,G14987,G14988,G14989,G14990,G14991,G14992,G14993,G14994,G14995,G14996,G14997,G14998,G14999,G15000,
       G15001,G15002,G15003,G15004,G15005,G15006,G15007,G15008,G15009,G15010,G15011,G15012,G15013,G15014,G15015,G15016,G15017,G15018,G15019,G15020,
       G15021,G15022,G15023,G15024,G15025,G15026,G15027,G15028,G15029,G15030,G15031,G15032,G15033,G15034,G15035,G15036,G15037,G15038,G15039,G15040,
       G15041,G15042,G15043,G15044,G15045,G15046,G15047,G15048,G15049,G15050,G15051,G15052,G15053,G15054,G15055,G15056,G15057,G15058,G15059,G15060,
       G15061,G15062,G15063,G15064,G15065,G15066,G15067,G15068,G15069,G15070,G15071,G15072,G15073,G15074,G15075,G15076,G15077,G15078,G15079,G15080,
       G15081,G15082,G15083,G15084,G15085,G15086,G15087,G15088,G15089,G15090,G15091,G15092,G15093,G15094,G15095,G15096,G15097,G15098,G15099,G15100,
       G15101,G15102,G15103,G15104,G15105,G15106,G15107,G15108,G15109,G15110,G15111,G15112,G15113,G15114,G15115,G15116,G15117,G15118,G15119,G15120,
       G15121,G15122,G15123,G15124,G15125,G15126,G15127,G15128,G15129,G15130,G15131,G15132,G15133,G15134,G15135,G15136,G15137,G15138,G15139,G15140,
       G15141,G15142,G15143,G15144,G15145,G15146,G15147,G15148,G15149,G15150,G15151,G15152,G15153,G15154,G15155,G15156,G15157,G15158,G15159,G15160,
       G15161,G15162,G15163,G15164,G15165,G15166,G15167,G15168,G15169,G15170,G15171,G15172,G15173,G15174,G15175,G15176,G15177,G15178,G15179,G15180,
       G15181,G15182,G15183,G15184,G15185,G15186,G15187,G15188,G15189,G15190,G15191,G15192,G15193,G15194,G15195,G15196,G15197,G15198,G15199,G15200,
       G15201,G15202,G15203,G15204,G15205,G15206,G15207,G15208,G15209,G15210,G15211,G15212,G15213,G15214,G15215,G15216,G15217,G15218,G15219,G15220,
       G15221,G15222,G15223,G15224,G15225,G15226,G15227,G15228,G15229,G15230,G15231,G15232,G15233,G15234,G15235,G15236,G15237,G15238,G15239,G15240,
       G15241,G15242,G15243,G15244,G15245,G15246,G15247,G15248,G15249,G15250,G15251,G15252,G15253,G15254,G15255,G15256,G15257,G15258,G15259,G15260,
       G15261,G15262,G15263,G15264,G15265,G15266,G15267,G15268,G15269,G15270,G15271,G15272,G15273,G15274,G15275,G15276,G15277,G15278,G15279,G15280,
       G15281,G15282,G15283,G15284,G15285,G15286,G15287,G15288,G15289,G15290,G15291,G15292,G15293,G15294,G15295,G15296,G15297,G15298,G15299,G15300,
       G15301,G15302,G15303,G15304,G15305,G15306,G15307,G15308,G15309,G15310,G15311,G15312,G15313,G15314,G15315,G15316,G15317,G15318,G15319,G15320,
       G15321,G15322,G15323,G15324,G15325,G15326,G15327,G15328,G15329,G15330,G15331,G15332,G15333,G15334,G15335,G15336,G15337,G15338,G15339,G15340,
       G15341,G15342,G15343,G15344,G15345,G15346,G15347,G15348,G15349,G15350,G15351,G15352,G15353,G15354,G15355,G15356,G15357,G15358,G15359,G15360,
       G15361,G15362,G15363,G15364,G15365,G15366,G15367,G15368,G15369,G15370,G15371,G15372,G15373,G15374,G15375,G15376,G15377,G15378,G15379,G15380,
       G15381,G15382,G15383,G15384,G15385,G15386,G15387,G15388,G15389,G15390,G15391,G15392,G15393,G15394,G15395,G15396,G15397,G15398,G15399,G15400,
       G15401,G15402,G15403,G15404,G15405,G15406,G15407,G15408,G15409,G15410,G15411,G15412,G15413,G15414,G15415,G15416,G15417,G15418,G15419,G15420,
       G15421,G15422,G15423,G15424,G15425,G15426,G15427,G15428,G15429,G15430,G15431,G15432,G15433,G15434,G15435,G15436,G15437,G15438,G15439,G15440,
       G15441,G15442,G15443,G15444,G15445,G15446,G15447,G15448,G15449,G15450,G15451,G15452,G15453,G15454,G15455,G15456,G15457,G15458,G15459,G15460,
       G15461,G15462,G15463,G15464,G15465,G15466,G15467,G15468,G15469,G15470,G15471,G15472,G15473,G15474,G15475,G15476,G15477,G15478,G15479,G15480,
       G15481,G15482,G15483,G15484,G15485,G15486,G15487,G15488,G15489,G15490,G15491,G15492,G15493,G15494,G15495,G15496,G15497,G15498,G15499,G15500,
       G15501,G15502,G15503,G15504,G15505,G15506,G15507,G15508,G15509,G15510,G15511,G15512,G15513,G15514,G15515,G15516,G15517,G15518,G15519,G15520,
       G15521,G15522,G15523,G15524,G15525,G15526,G15527,G15528,G15529,G15530,G15531,G15532,G15533,G15534,G15535,G15536,G15537,G15538,G15539,G15540,
       G15541,G15542,G15543,G15544,G15545,G15546,G15547,G15548,G15549,G15550,G15551,G15552,G15553,G15554,G15555,G15556,G15557,G15558,G15559,G15560,
       G15561,G15562,G15563,G15564,G15565,G15566,G15567,G15568,G15569,G15570,G15571,G15572,G15573,G15574,G15575,G15576,G15577,G15578,G15579,G15580,
       G15581,G15582,G15583,G15584,G15585,G15586,G15587,G15588,G15589,G15590,G15591,G15592,G15593,G15594,G15595,G15596,G15597,G15598,G15599,G15600,
       G15601,G15602,G15603,G15604,G15605,G15606,G15607,G15608,G15609,G15610,G15611,G15612,G15613,G15614,G15615,G15616,G15617,G15618,G15619,G15620,
       G15621,G15622,G15623,G15624,G15625,G15626,G15627,G15628,G15629,G15630,G15631,G15632,G15633,G15634,G15635,G15636,G15637,G15638,G15639,G15640,
       G15641,G15642,G15643,G15644,G15645,G15646,G15647,G15648,G15649,G15650,G15651,G15652,G15653,G15654,G15655,G15656,G15657,G15658,G15659,G15660,
       G15661,G15662,G15663,G15664,G15665,G15666,G15667,G15668,G15669,G15670,G15671,G15672,G15673,G15674,G15675,G15676,G15677,G15678,G15679,G15680,
       G15681,G15682,G15683,G15684,G15685,G15686,G15687,G15688,G15689,G15690,G15691,G15692,G15693,G15694,G15695,G15696,G15697,G15698,G15699,G15700,
       G15701,G15702,G15703,G15704,G15705,G15706,G15707,G15708,G15709,G15710,G15711,G15712,G15713,G15714,G15715,G15716,G15717,G15718,G15719,G15720,
       G15721,G15722,G15723,G15724,G15725,G15726,G15727,G15728,G15729,G15730,G15731,G15732,G15733,G15734,G15735,G15736,G15737,G15738,G15739,G15740,
       G15741,G15742,G15743,G15744,G15745,G15746,G15747,G15748,G15749,G15750,G15751,G15752,G15753,G15754,G15755,G15756,G15757,G15758,G15759,G15760,
       G15761,G15762,G15763,G15764,G15765,G15766,G15767,G15768,G15769,G15770,G15771,G15772,G15773,G15774,G15775,G15776,G15777,G15778,G15779,G15780,
       G15781,G15782,G15783,G15784,G15785,G15786,G15787,G15788,G15789,G15790,G15791,G15792,G15793,G15794,G15795,G15796,G15797,G15798,G15799,G15800,
       G15801,G15802,G15803,G15804,G15805,G15806,G15807,G15808,G15809,G15810,G15811,G15812,G15813,G15814,G15815,G15816,G15817,G15818,G15819,G15820,
       G15821,G15822,G15823,G15824,G15825,G15826,G15827,G15828,G15829,G15830,G15831,G15832,G15833,G15834,G15835,G15836,G15837,G15838,G15839,G15840,
       G15841,G15842,G15843,G15844,G15845,G15846,G15847,G15848,G15849,G15850,G15851,G15852,G15853,G15854,G15855,G15856,G15857,G15858,G15859,G15860,
       G15861,G15862,G15863,G15864,G15865,G15866,G15867,G15868,G15869,G15870,G15871,G15872,G15873,G15874,G15875,G15876,G15877,G15878,G15879,G15880,
       G15881,G15882,G15883,G15884,G15885,G15886,G15887,G15888,G15889,G15890,G15891,G15892,G15893,G15894,G15895,G15896,G15897,G15898,G15899,G15900,
       G15901,G15902,G15903,G15904,G15905,G15906,G15907,G15908,G15909,G15910,G15911,G15912,G15913,G15914,G15915,G15916,G15917,G15918,G15919,G15920,
       G15921,G15922,G15923,G15924,G15925,G15926,G15927,G15928,G15929,G15930,G15931,G15932,G15933,G15934,G15935,G15936,G15937,G15938,G15939,G15940,
       G15941,G15942,G15943,G15944,G15945,G15946,G15947,G15948,G15949,G15950,G15951,G15952,G15953,G15954,G15955,G15956,G15957,G15958,G15959,G15960,
       G15961,G15962,G15963,G15964,G15965,G15966,G15967,G15968,G15969,G15970,G15971,G15972,G15973,G15974,G15975,G15976,G15977,G15978,G15979,G15980,
       G15981,G15982,G15983,G15984,G15985,G15986,G15987,G15988,G15989,G15990,G15991,G15992,G15993,G15994,G15995,G15996,G15997,G15998,G15999,G16000,
       G16001,G16002,G16003,G16004,G16005,G16006,G16007,G16008,G16009,G16010,G16011,G16012,G16013,G16014,G16015,G16016,G16017,G16018,G16019,G16020,
       G16021,G16022,G16023,G16024,G16025,G16026,G16027,G16028,G16029,G16030,G16031,G16032,G16033,G16034,G16035,G16036,G16037,G16038,G16039,G16040,
       G16041,G16042,G16043,G16044,G16045,G16046,G16047,G16048,G16049,G16050,G16051,G16052,G16053,G16054,G16055,G16056,G16057,G16058,G16059,G16060,
       G16061,G16062,G16063,G16064,G16065,G16066,G16067,G16068,G16069,G16070,G16071,G16072,G16073,G16074,G16075,G16076,G16077,G16078,G16079,G16080,
       G16081,G16082,G16083,G16084,G16085,G16086,G16087,G16088,G16089,G16090,G16091,G16092,G16093,G16094,G16095,G16096,G16097,G16098,G16099,G16100,
       G16101,G16102,G16103,G16104,G16105,G16106,G16107,G16108,G16109,G16110,G16111,G16112,G16113,G16114,G16115,G16116,G16117,G16118,G16119,G16120,
       G16121,G16122,G16123,G16124,G16125,G16126,G16127,G16128,G16129,G16130,G16131,G16132,G16133,G16134,G16135,G16136,G16137,G16138,G16139,G16140,
       G16141,G16142,G16143,G16144,G16145,G16146,G16147,G16148,G16149,G16150,G16151,G16152,G16153,G16154,G16155,G16156,G16157,G16158,G16159,G16160,
       G16161,G16162,G16163,G16164,G16165,G16166,G16167,G16168,G16169,G16170,G16171,G16172,G16173,G16174,G16175,G16176,G16177,G16178,G16179,G16180,
       G16181,G16182,G16183,G16184,G16185,G16186,G16187,G16188,G16189,G16190,G16191,G16192,G16193,G16194,G16195,G16196,G16197,G16198,G16199,G16200,
       G16201,G16202,G16203,G16204,G16205,G16206,G16207,G16208,G16209,G16210,G16211,G16212,G16213,G16214,G16215,G16216,G16217,G16218,G16219,G16220,
       G16221,G16222,G16223,G16224,G16225,G16226,G16227,G16228,G16229,G16230,G16231,G16232,G16233,G16234,G16235,G16236,G16237,G16238,G16239,G16240,
       G16241,G16242,G16243,G16244,G16245,G16246,G16247,G16248,G16249,G16250,G16251,G16252,G16253,G16254,G16255,G16256,G16257,G16258,G16259,G16260,
       G16261,G16262,G16263,G16264,G16265,G16266,G16267,G16268,G16269,G16270,G16271,G16272,G16273,G16274,G16275,G16276,G16277,G16278,G16279,G16280,
       G16281,G16282,G16283,G16284,G16285,G16286,G16287,G16288,G16289,G16290,G16291,G16292,G16293,G16294,G16295,G16296,G16297,G16298,G16299,G16300,
       G16301,G16302,G16303,G16304,G16305,G16306,G16307,G16308,G16309,G16310,G16311,G16312,G16313,G16314,G16315,G16316,G16317,G16318,G16319,G16320,
       G16321,G16322,G16323,G16324,G16325,G16326,G16327,G16328,G16329,G16330,G16331,G16332,G16333,G16334,G16335,G16336,G16337,G16338,G16339,G16340,
       G16341,G16342,G16343,G16344,G16345,G16346,G16347,G16348,G16349,G16350,G16351,G16352,G16353,G16354,G16355,G16356,G16357,G16358,G16359,G16360,
       G16361,G16362,G16363,G16364,G16365,G16366,G16367,G16368,G16369,G16370,G16371,G16372,G16373,G16374,G16375,G16376,G16377,G16378,G16379,G16380,
       G16381,G16382,G16383,G16384,G16385,G16386,G16387,G16388,G16389,G16390,G16391,G16392,G16393,G16394,G16395,G16396,G16397,G16398,G16399,G16400,
       G16401,G16402,G16403,G16404,G16405,G16406,G16407,G16408,G16409,G16410,G16411,G16412,G16413,G16414,G16415,G16416,G16417,G16418,G16419,G16420,
       G16421,G16422,G16423,G16424,G16425,G16426,G16427,G16428,G16429,G16430,G16431,G16432,G16433,G16434,G16435,G16436,G16437,G16438,G16439,G16440,
       G16441,G16442,G16443,G16444,G16445,G16446,G16447,G16448,G16449,G16450,G16451,G16452,G16453,G16454,G16455,G16456,G16457,G16458,G16459,G16460,
       G16461,G16462,G16463,G16464,G16465,G16466,G16467,G16468,G16469,G16470,G16471,G16472,G16473,G16474,G16475,G16476,G16477,G16478,G16479,G16480,
       G16481,G16482,G16483,G16484,G16485,G16486,G16487,G16488,G16489,G16490,G16491,G16492,G16493,G16494,G16495,G16496,G16497,G16498,G16499,G16500,
       G16501,G16502,G16503,G16504,G16505,G16506,G16507,G16508,G16509,G16510,G16511,G16512,G16513,G16514,G16515,G16516,G16517,G16518,G16519,G16520,
       G16521,G16522,G16523,G16524,G16525,G16526,G16527,G16528,G16529,G16530,G16531,G16532,G16533,G16534,G16535,G16536,G16537,G16538,G16539,G16540,
       G16541,G16542,G16543,G16544,G16545,G16546,G16547,G16548,G16549,G16550,G16551,G16552,G16553,G16554,G16555,G16556,G16557,G16558,G16559,G16560,
       G16561,G16562,G16563,G16564,G16565,G16566,G16567,G16568,G16569,G16570,G16571,G16572,G16573,G16574,G16575,G16576,G16577,G16578,G16579,G16580,
       G16581,G16582,G16583,G16584,G16585,G16586,G16587,G16588,G16589,G16590,G16591,G16592,G16593,G16594,G16595,G16596,G16597,G16598,G16599,G16600,
       G16601,G16602,G16603,G16604,G16605,G16606,G16607,G16608,G16609,G16610,G16611,G16612,G16613,G16614,G16615,G16616,G16617,G16618,G16619,G16620,
       G16621,G16622,G16623,G16624,G16625,G16626,G16627,G16628,G16629,G16630,G16631,G16632,G16633,G16634,G16635,G16636,G16637,G16638,G16639,G16640,
       G16641,G16642,G16643,G16644,G16645,G16646,G16647,G16648,G16649,G16650,G16651,G16652,G16653,G16654,G16655,G16656,G16657,G16658,G16659,G16660,
       G16661,G16662,G16663,G16664,G16665,G16666,G16667,G16668,G16669,G16670,G16671,G16672,G16673,G16674,G16675,G16676,G16677,G16678,G16679,G16680,
       G16681,G16682,G16683,G16684,G16685,G16686,G16687,G16688,G16689,G16690,G16691,G16692,G16693,G16694,G16695,G16696,G16697,G16698,G16699,G16700,
       G16701,G16702,G16703,G16704,G16705,G16706,G16707,G16708,G16709,G16710,G16711,G16712,G16713,G16714,G16715,G16716,G16717,G16718,G16719,G16720,
       G16721,G16722,G16723,G16724,G16725,G16726,G16727,G16728,G16729,G16730,G16731,G16732,G16733,G16734,G16735,G16736,G16737,G16738,G16739,G16740,
       G16741,G16742,G16743,G16744,G16745,G16746,G16747,G16748,G16749,G16750,G16751,G16752,G16753,G16754,G16755,G16756,G16757,G16758,G16759,G16760,
       G16761,G16762,G16763,G16764,G16765,G16766,G16767,G16768,G16769,G16770,G16771,G16772,G16773,G16774,G16775,G16776,G16777,G16778,G16779,G16780,
       G16781,G16782,G16783,G16784,G16785,G16786,G16787,G16788,G16789,G16790,G16791,G16792,G16793,G16794,G16795,G16796,G16797,G16798,G16799,G16800,
       G16801,G16802,G16803,G16804,G16805,G16806,G16807,G16808,G16809,G16810,G16811,G16812,G16813,G16814,G16815,G16816,G16817,G16818,G16819,G16820,
       G16821,G16822,G16823,G16824,G16825,G16826,G16827,G16828,G16829,G16830,G16831,G16832,G16833,G16834,G16835,G16836,G16837,G16838,G16839,G16840,
       G16841,G16842,G16843,G16844,G16845,G16846,G16847,G16848,G16849,G16850,G16851,G16852,G16853,G16854,G16855,G16856,G16857,G16858,G16859,G16860,
       G16861,G16862,G16863,G16864,G16865,G16866,G16867,G16868,G16869,G16870,G16871,G16872,G16873,G16874,G16875,G16876,G16877,G16878,G16879,G16880,
       G16881,G16882,G16883,G16884,G16885,G16886,G16887,G16888,G16889,G16890,G16891,G16892,G16893,G16894,G16895,G16896,G16897,G16898,G16899,G16900,
       G16901,G16902,G16903,G16904,G16905,G16906,G16907,G16908,G16909,G16910,G16911,G16912,G16913,G16914,G16915,G16916,G16917,G16918,G16919,G16920,
       G16921,G16922,G16923,G16924,G16925,G16926,G16927,G16928,G16929,G16930,G16931,G16932,G16933,G16934,G16935,G16936,G16937,G16938,G16939,G16940,
       G16941,G16942,G16943,G16944,G16945,G16946,G16947,G16948,G16949,G16950,G16951,G16952,G16953,G16954,G16955,G16956,G16957,G16958,G16959,G16960,
       G16961,G16962,G16963,G16964,G16965,G16966,G16967,G16968,G16969,G16970,G16971,G16972,G16973,G16974,G16975,G16976,G16977,G16978,G16979,G16980,
       G16981,G16982,G16983,G16984,G16985,G16986,G16987,G16988,G16989,G16990,G16991,G16992,G16993,G16994,G16995,G16996,G16997,G16998,G16999,G17000,
       G17001,G17002,G17003,G17004,G17005,G17006,G17007,G17008,G17009,G17010,G17011,G17012,G17013,G17014,G17015,G17016,G17017,G17018,G17019,G17020,
       G17021,G17022,G17023,G17024,G17025,G17026,G17027,G17028,G17029,G17030,G17031,G17032,G17033,G17034,G17035,G17036,G17037,G17038,G17039,G17040,
       G17041,G17042,G17043,G17044,G17045,G17046,G17047,G17048,G17049,G17050,G17051,G17052,G17053,G17054,G17055,G17056,G17057,G17058,G17059,G17060,
       G17061,G17062,G17063,G17064,G17065,G17066,G17067,G17068,G17069,G17070,G17071,G17072,G17073,G17074,G17075,G17076,G17077,G17078,G17079,G17080,
       G17081,G17082,G17083,G17084,G17085,G17086,G17087,G17088,G17089,G17090,G17091,G17092,G17093,G17094,G17095,G17096,G17097,G17098,G17099,G17100,
       G17101,G17102,G17103,G17104,G17105,G17106,G17107,G17108,G17109,G17110,G17111,G17112,G17113,G17114,G17115,G17116,G17117,G17118,G17119,G17120,
       G17121,G17122,G17123,G17124,G17125,G17126,G17127,G17128,G17129,G17130,G17131,G17132,G17133,G17134,G17135,G17136,G17137,G17138,G17139,G17140,
       G17141,G17142,G17143,G17144,G17145,G17146,G17147,G17148,G17149,G17150,G17151,G17152,G17153,G17154,G17155,G17156,G17157,G17158,G17159,G17160,
       G17161,G17162,G17163,G17164,G17165,G17166,G17167,G17168,G17169,G17170,G17171,G17172,G17173,G17174,G17175,G17176,G17177,G17178,G17179,G17180,
       G17181,G17182,G17183,G17184,G17185,G17186,G17187,G17188,G17189,G17190,G17191,G17192,G17193,G17194,G17195,G17196,G17197,G17198,G17199,G17200,
       G17201,G17202,G17203,G17204,G17205,G17206,G17207,G17208,G17209,G17210,G17211,G17212,G17213,G17214,G17215,G17216,G17217,G17218,G17219,G17220,
       G17221,G17222,G17223,G17224,G17225,G17226,G17227,G17228,G17229,G17230,G17231,G17232,G17233,G17234,G17235,G17236,G17237,G17238,G17239,G17240,
       G17241,G17242,G17243,G17244,G17245,G17246,G17247,G17248,G17249,G17250,G17251,G17252,G17253,G17254,G17255,G17256,G17257,G17258,G17259,G17260,
       G17261,G17262,G17263,G17264,G17265,G17266,G17267,G17268,G17269,G17270,G17271,G17272,G17273,G17274,G17275,G17276,G17277,G17278,G17279,G17280,
       G17281,G17282,G17283,G17284,G17285,G17286,G17287,G17288,G17289,G17290,G17291,G17292,G17293,G17294,G17295,G17296,G17297,G17298,G17299,G17300,
       G17301,G17302,G17303,G17304,G17305,G17306,G17307,G17308,G17309,G17310,G17311,G17312,G17313,G17314,G17315,G17316,G17317,G17318,G17319,G17320,
       G17321,G17322,G17323,G17324,G17325,G17326,G17327,G17328,G17329,G17330,G17331,G17332,G17333,G17334,G17335,G17336,G17337,G17338,G17339,G17340,
       G17341,G17342,G17343,G17344,G17345,G17346,G17347,G17348,G17349,G17350,G17351,G17352,G17353,G17354,G17355,G17356,G17357,G17358,G17359,G17360,
       G17361,G17362,G17363,G17364,G17365,G17366,G17367,G17368,G17369,G17370,G17371,G17372,G17373,G17374,G17375,G17376,G17377,G17378,G17379,G17380,
       G17381,G17382,G17383,G17384,G17385,G17386,G17387,G17388,G17389,G17390,G17391,G17392,G17393,G17394,G17395,G17396,G17397,G17398,G17399,G17400,
       G17401,G17402,G17403,G17404,G17405,G17406,G17407,G17408,G17409,G17410,G17411,G17412,G17413,G17414,G17415,G17416,G17417,G17418,G17419,G17420,
       G17421,G17422,G17423,G17424,G17425,G17426,G17427,G17428,G17429,G17430,G17431,G17432,G17433,G17434,G17435,G17436,G17437,G17438,G17439,G17440,
       G17441,G17442,G17443,G17444,G17445,G17446,G17447,G17448,G17449,G17450,G17451,G17452,G17453,G17454,G17455,G17456,G17457,G17458,G17459,G17460,
       G17461,G17462,G17463,G17464,G17465,G17466,G17467,G17468,G17469,G17470,G17471,G17472,G17473,G17474,G17475,G17476,G17477,G17478,G17479,G17480,
       G17481,G17482,G17483,G17484,G17485,G17486,G17487,G17488,G17489,G17490,G17491,G17492,G17493,G17494,G17495,G17496,G17497,G17498,G17499,G17500,
       G17501,G17502,G17503,G17504,G17505,G17506,G17507,G17508,G17509,G17510,G17511,G17512,G17513,G17514,G17515,G17516,G17517,G17518,G17519,G17520,
       G17521,G17522,G17523,G17524,G17525,G17526,G17527,G17528,G17529,G17530,G17531,G17532,G17533,G17534,G17535,G17536,G17537,G17538,G17539,G17540,
       G17541,G17542,G17543,G17544,G17545,G17546,G17547,G17548,G17549,G17550,G17551,G17552,G17553,G17554,G17555,G17556,G17557,G17558,G17559,G17560,
       G17561,G17562,G17563,G17564,G17565,G17566,G17567,G17568,G17569,G17570,G17571,G17572,G17573,G17574,G17575,G17576,G17577,G17578,G17579,G17580,
       G17581,G17582,G17583,G17584,G17585,G17586,G17587,G17588,G17589,G17590,G17591,G17592,G17593,G17594,G17595,G17596,G17597,G17598,G17599,G17600,
       G17601,G17602,G17603,G17604,G17605,G17606,G17607,G17608,G17609,G17610,G17611,G17612,G17613,G17614,G17615,G17616,G17617,G17618,G17619,G17620,
       G17621,G17622,G17623,G17624,G17625,G17626,G17627,G17628,G17629,G17630,G17631,G17632,G17633,G17634,G17635,G17636,G17637,G17638,G17639,G17640,
       G17641,G17642,G17643,G17644,G17645,G17646,G17647,G17648,G17649,G17650,G17651,G17652,G17653,G17654,G17655,G17656,G17657,G17658,G17659,G17660,
       G17661,G17662,G17663,G17664,G17665,G17666,G17667,G17668,G17669,G17670,G17671,G17672,G17673,G17674,G17675,G17676,G17677,G17678,G17679,G17680,
       G17681,G17682,G17683,G17684,G17685,G17686,G17687,G17688,G17689,G17690,G17691,G17692,G17693,G17694,G17695,G17696,G17697,G17698,G17699,G17700,
       G17701,G17702,G17703,G17704,G17705,G17706,G17707,G17708,G17709,G17710,G17711,G17712,G17713,G17714,G17715,G17716,G17717,G17718,G17719,G17720,
       G17721,G17722,G17723,G17724,G17725,G17726,G17727,G17728,G17729,G17730,G17731,G17732,G17733,G17734,G17735,G17736,G17737,G17738,G17739,G17740,
       G17741,G17742,G17743,G17744,G17745,G17746,G17747,G17748,G17749,G17750,G17751,G17752,G17753,G17754,G17755,G17756,G17757,G17758,G17759,G17760,
       G17761,G17762,G17763,G17764,G17765,G17766,G17767,G17768,G17769,G17770,G17771,G17772,G17773,G17774,G17775,G17776,G17777,G17778,G17779,G17780,
       G17781,G17782,G17783,G17784,G17785,G17786,G17787,G17788,G17789,G17790,G17791,G17792,G17793,G17794,G17795,G17796,G17797,G17798,G17799,G17800,
       G17801,G17802,G17803,G17804,G17805,G17806,G17807,G17808,G17809,G17810,G17811,G17812,G17813,G17814,G17815,G17816,G17817,G17818,G17819,G17820,
       G17821,G17822,G17823,G17824,G17825,G17826,G17827,G17828,G17829,G17830,G17831,G17832,G17833,G17834,G17835,G17836,G17837,G17838,G17839,G17840,
       G17841,G17842,G17843,G17844,G17845,G17846,G17847,G17848,G17849,G17850,G17851,G17852,G17853,G17854,G17855,G17856,G17857,G17858,G17859,G17860,
       G17861,G17862,G17863,G17864,G17865,G17866,G17867,G17868,G17869,G17870,G17871,G17872,G17873,G17874,G17875,G17876,G17877,G17878,G17879,G17880,
       G17881,G17882,G17883,G17884,G17885,G17886,G17887,G17888,G17889,G17890,G17891,G17892,G17893,G17894,G17895,G17896,G17897,G17898,G17899,G17900,
       G17901,G17902,G17903,G17904,G17905,G17906,G17907,G17908,G17909,G17910,G17911,G17912,G17913,G17914,G17915,G17916,G17917,G17918,G17919,G17920,
       G17921,G17922,G17923,G17924,G17925,G17926,G17927,G17928,G17929,G17930,G17931,G17932,G17933,G17934,G17935,G17936,G17937,G17938,G17939,G17940,
       G17941,G17942,G17943,G17944,G17945,G17946,G17947,G17948,G17949,G17950,G17951,G17952,G17953,G17954,G17955,G17956,G17957,G17958,G17959,G17960,
       G17961,G17962,G17963,G17964,G17965,G17966,G17967,G17968,G17969,G17970,G17971,G17972,G17973,G17974,G17975,G17976,G17977,G17978,G17979,G17980,
       G17981,G17982,G17983,G17984,G17985,G17986,G17987,G17988,G17989,G17990,G17991,G17992,G17993,G17994,G17995,G17996,G17997,G17998,G17999,G18000,
       G18001,G18002,G18003,G18004,G18005,G18006,G18007,G18008,G18009,G18010,G18011,G18012,G18013,G18014,G18015,G18016,G18017,G18018,G18019,G18020,
       G18021,G18022,G18023,G18024,G18025,G18026,G18027,G18028,G18029,G18030,G18031,G18032,G18033,G18034,G18035,G18036,G18037,G18038,G18039,G18040,
       G18041,G18042,G18043,G18044,G18045,G18046,G18047,G18048,G18049,G18050,G18051,G18052,G18053,G18054,G18055,G18056,G18057,G18058,G18059,G18060,
       G18061,G18062,G18063,G18064,G18065,G18066,G18067,G18068,G18069,G18070,G18071,G18072,G18073,G18074,G18075,G18076,G18077,G18078,G18079,G18080,
       G18081,G18082,G18083,G18084,G18085,G18086,G18087,G18088,G18089,G18090,G18091,G18092,G18093,G18094,G18095,G18096,G18097,G18098,G18099,G18100,
       G18101,G18102,G18103,G18104,G18105,G18106,G18107,G18108,G18109,G18110,G18111,G18112,G18113,G18114,G18115,G18116,G18117,G18118,G18119,G18120,
       G18121,G18122,G18123,G18124,G18125,G18126,G18127,G18128,G18129,G18130,G18131,G18132,G18133,G18134,G18135,G18136,G18137,G18138,G18139,G18140,
       G18141,G18142,G18143,G18144,G18145,G18146,G18147,G18148,G18149,G18150,G18151,G18152,G18153,G18154,G18155,G18156,G18157,G18158,G18159,G18160,
       G18161,G18162,G18163,G18164,G18165,G18166,G18167,G18168,G18169,G18170,G18171,G18172,G18173,G18174,G18175,G18176,G18177,G18178,G18179,G18180,
       G18181,G18182,G18183,G18184,G18185,G18186,G18187,G18188,G18189,G18190,G18191,G18192,G18193,G18194,G18195,G18196,G18197,G18198,G18199,G18200,
       G18201,G18202,G18203,G18204,G18205,G18206,G18207,G18208,G18209,G18210,G18211,G18212,G18213,G18214,G18215,G18216,G18217,G18218,G18219,G18220,
       G18221,G18222,G18223,G18224,G18225,G18226,G18227,G18228,G18229,G18230,G18231,G18232,G18233,G18234,G18235,G18236,G18237,G18238,G18239,G18240,
       G18241,G18242,G18243,G18244,G18245,G18246,G18247,G18248,G18249,G18250,G18251,G18252,G18253,G18254,G18255,G18256,G18257,G18258,G18259,G18260,
       G18261,G18262,G18263,G18264,G18265,G18266,G18267,G18268,G18269,G18270,G18271,G18272,G18273,G18274,G18275,G18276,G18277,G18278,G18279,G18280,
       G18281,G18282,G18283,G18284,G18285,G18286,G18287,G18288,G18289,G18290,G18291,G18292,G18293,G18294,G18295,G18296,G18297,G18298,G18299,G18300,
       G18301,G18302,G18303,G18304,G18305,G18306,G18307,G18308,G18309,G18310,G18311,G18312,G18313,G18314,G18315,G18316,G18317,G18318,G18319,G18320,
       G18321,G18322,G18323,G18324,G18325,G18326,G18327,G18328,G18329,G18330,G18331,G18332,G18333,G18334,G18335,G18336,G18337,G18338,G18339,G18340,
       G18341,G18342,G18343,G18344,G18345,G18346,G18347,G18348,G18349,G18350,G18351,G18352,G18353,G18354,G18355,G18356,G18357,G18358,G18359,G18360,
       G18361,G18362,G18363,G18364,G18365,G18366,G18367,G18368,G18369,G18370,G18371,G18372,G18373,G18374,G18375,G18376,G18377,G18378,G18379,G18380,
       G18381,G18382,G18383,G18384,G18385,G18386,G18387,G18388,G18389,G18390,G18391,G18392,G18393,G18394,G18395,G18396,G18397,G18398,G18399,G18400,
       G18401,G18402,G18403,G18404,G18405,G18406,G18407,G18408,G18409,G18410,G18411,G18412,G18413,G18414,G18415,G18416,G18417,G18418,G18419,G18420,
       G18421,G18422,G18423,G18424,G18425,G18426,G18427,G18428,G18429,G18430,G18431,G18432,G18433,G18434,G18435,G18436,G18437,G18438,G18439,G18440,
       G18441,G18442,G18443,G18444,G18445,G18446,G18447,G18448,G18449,G18450,G18451,G18452,G18453,G18454,G18455,G18456,G18457,G18458,G18459,G18460,
       G18461,G18462,G18463,G18464,G18465,G18466,G18467,G18468,G18469,G18470,G18471,G18472,G18473,G18474,G18475,G18476,G18477,G18478,G18479,G18480,
       G18481,G18482,G18483,G18484,G18485,G18486,G18487,G18488,G18489,G18490,G18491,G18492,G18493,G18494,G18495,G18496,G18497,G18498,G18499,G18500,
       G18501,G18502,G18503,G18504,G18505,G18506,G18507,G18508,G18509,G18510,G18511,G18512,G18513,G18514,G18515,G18516,G18517,G18518,G18519,G18520,
       G18521,G18522,G18523,G18524,G18525,G18526,G18527,G18528,G18529,G18530,G18531,G18532,G18533,G18534,G18535,G18536,G18537,G18538,G18539,G18540,
       G18541,G18542,G18543,G18544,G18545,G18546,G18547,G18548,G18549,G18550,G18551,G18552,G18553,G18554,G18555,G18556,G18557,G18558,G18559,G18560,
       G18561,G18562,G18563,G18564,G18565,G18566,G18567,G18568,G18569,G18570,G18571,G18572,G18573,G18574,G18575,G18576,G18577,G18578,G18579,G18580,
       G18581,G18582,G18583,G18584,G18585,G18586,G18587,G18588,G18589,G18590,G18591,G18592,G18593,G18594,G18595,G18596,G18597,G18598,G18599,G18600,
       G18601,G18602,G18603,G18604,G18605,G18606,G18607,G18608,G18609,G18610,G18611,G18612,G18613,G18614,G18615,G18616,G18617,G18618,G18619,G18620,
       G18621,G18622,G18623,G18624,G18625,G18626,G18627,G18628,G18629,G18630,G18631,G18632,G18633,G18634,G18635,G18636,G18637,G18638,G18639,G18640,
       G18641,G18642,G18643,G18644,G18645,G18646,G18647,G18648,G18649,G18650,G18651,G18652,G18653,G18654,G18655,G18656,G18657,G18658,G18659,G18660,
       G18661,G18662,G18663,G18664,G18665,G18666,G18667,G18668,G18669,G18670,G18671,G18672,G18673,G18674,G18675,G18676,G18677,G18678,G18679,G18680,
       G18681,G18682,G18683,G18684,G18685,G18686,G18687,G18688,G18689,G18690,G18691,G18692,G18693,G18694,G18695,G18696,G18697,G18698,G18699,G18700,
       G18701,G18702,G18703,G18704,G18705,G18706,G18707,G18708,G18709,G18710,G18711,G18712,G18713,G18714,G18715,G18716,G18717,G18718,G18719,G18720,
       G18721,G18722,G18723,G18724,G18725,G18726,G18727,G18728,G18729,G18730,G18731,G18732,G18733,G18734,G18735,G18736,G18737,G18738,G18739,G18740,
       G18741,G18742,G18743,G18744,G18745,G18746,G18747,G18748,G18749,G18750,G18751,G18752,G18753,G18754,G18755,G18756,G18757,G18758,G18759,G18760,
       G18761,G18762,G18763,G18764,G18765,G18766,G18767,G18768,G18769,G18770,G18771,G18772,G18773,G18774,G18775,G18776,G18777,G18778,G18779,G18780,
       G18781,G18782,G18783,G18784,G18785,G18786,G18787,G18788,G18789,G18790,G18791,G18792,G18793,G18794,G18795,G18796,G18797,G18798,G18799,G18800,
       G18801,G18802,G18803,G18804,G18805,G18806,G18807,G18808,G18809,G18810,G18811,G18812,G18813,G18814,G18815,G18816,G18817,G18818,G18819,G18820,
       G18821,G18822,G18823,G18824,G18825,G18826,G18827,G18828,G18829,G18830,G18831,G18832,G18833,G18834,G18835,G18836,G18837,G18838,G18839,G18840,
       G18841,G18842,G18843,G18844,G18845,G18846,G18847,G18848,G18849,G18850,G18851,G18852,G18853,G18854,G18855,G18856,G18857,G18858,G18859,G18860,
       G18861,G18862,G18863,G18864,G18865,G18866,G18867,G18868,G18869,G18870,G18871,G18872,G18873,G18874,G18875,G18876,G18877,G18878,G18879,G18880,
       G18881,G18882,G18883,G18884,G18885,G18886,G18887,G18888,G18889,G18890,G18891,G18892,G18893,G18894,G18895,G18896,G18897,G18898,G18899,G18900,
       G18901,G18902,G18903,G18904,G18905,G18906,G18907,G18908,G18909,G18910,G18911,G18912,G18913,G18914,G18915,G18916,G18917,G18918,G18919,G18920,
       G18921,G18922,G18923,G18924,G18925,G18926,G18927,G18928,G18929,G18930,G18931,G18932,G18933,G18934,G18935,G18936,G18937,G18938,G18939,G18940,
       G18941,G18942,G18943,G18944,G18945,G18946,G18947,G18948,G18949,G18950,G18951,G18952,G18953,G18954,G18955,G18956,G18957,G18958,G18959,G18960,
       G18961,G18962,G18963,G18964,G18965,G18966,G18967,G18968,G18969,G18970,G18971,G18972,G18973,G18974,G18975,G18976,G18977,G18978,G18979,G18980,
       G18981,G18982,G18983,G18984,G18985,G18986,G18987,G18988,G18989,G18990,G18991,G18992,G18993,G18994,G18995,G18996,G18997,G18998,G18999,G19000,
       G19001,G19002,G19003,G19004,G19005,G19006,G19007,G19008,G19009,G19010,G19011,G19012,G19013,G19014,G19015,G19016,G19017,G19018,G19019,G19020,
       G19021,G19022,G19023,G19024,G19025,G19026,G19027,G19028,G19029,G19030,G19031,G19032,G19033,G19034,G19035,G19036,G19037,G19038,G19039,G19040,
       G19041,G19042,G19043,G19044,G19045,G19046,G19047,G19048,G19049,G19050,G19051,G19052,G19053,G19054,G19055,G19056,G19057,G19058,G19059,G19060,
       G19061,G19062,G19063,G19064,G19065,G19066,G19067,G19068,G19069,G19070,G19071,G19072,G19073,G19074,G19075,G19076,G19077,G19078,G19079,G19080,
       G19081,G19082,G19083,G19084,G19085,G19086,G19087,G19088,G19089,G19090,G19091,G19092,G19093,G19094,G19095,G19096,G19097,G19098,G19099,G19100,
       G19101,G19102,G19103,G19104,G19105,G19106,G19107,G19108,G19109,G19110,G19111,G19112,G19113,G19114,G19115,G19116,G19117,G19118,G19119,G19120,
       G19121,G19122,G19123,G19124,G19125,G19126,G19127,G19128,G19129,G19130,G19131,G19132,G19133,G19134,G19135,G19136,G19137,G19138,G19139,G19140,
       G19141,G19142,G19143,G19144,G19145,G19146,G19147,G19148,G19149,G19150,G19151,G19152,G19153,G19154,G19155,G19156,G19157,G19158,G19159,G19160,
       G19161,G19162,G19163,G19164,G19165,G19166,G19167,G19168,G19169,G19170,G19171,G19172,G19173,G19174,G19175,G19176,G19177,G19178,G19179,G19180,
       G19181,G19182,G19183,G19184,G19185,G19186,G19187,G19188,G19189,G19190,G19191,G19192,G19193,G19194,G19195,G19196,G19197,G19198,G19199,G19200,
       G19201,G19202,G19203,G19204,G19205,G19206,G19207,G19208,G19209,G19210,G19211,G19212,G19213,G19214,G19215,G19216,G19217,G19218,G19219,G19220,
       G19221,G19222,G19223,G19224,G19225,G19226,G19227,G19228,G19229,G19230,G19231,G19232,G19233,G19234,G19235,G19236,G19237,G19238,G19239,G19240,
       G19241,G19242,G19243,G19244,G19245,G19246,G19247,G19248,G19249,G19250,G19251,G19252,G19253,G19254,G19255,G19256,G19257,G19258,G19259,G19260,
       G19261,G19262,G19263,G19264,G19265,G19266,G19267,G19268,G19269,G19270,G19271,G19272,G19273,G19274,G19275,G19276,G19277,G19278,G19279,G19280,
       G19281,G19282,G19283,G19284,G19285,G19286,G19287,G19288,G19289,G19290,G19291,G19292,G19293,G19294,G19295,G19296,G19297,G19298,G19299,G19300,
       G19301,G19302,G19303,G19304,G19305,G19306,G19307,G19308,G19309,G19310,G19311,G19312,G19313,G19314,G19315,G19316,G19317,G19318,G19319,G19320,
       G19321,G19322,G19323,G19324,G19325,G19326,G19327,G19328,G19329,G19330,G19331,G19332,G19333,G19334,G19335,G19336,G19337,G19338,G19339,G19340,
       G19341,G19342,G19343,G19344,G19345,G19346,G19347,G19348,G19349,G19350,G19351,G19352,G19353,G19354,G19355,G19356,G19357,G19358,G19359,G19360,
       G19361,G19362,G19363,G19364,G19365,G19366,G19367,G19368,G19369,G19370,G19371,G19372,G19373,G19374,G19375,G19376,G19377,G19378,G19379,G19380,
       G19381,G19382,G19383,G19384,G19385,G19386,G19387,G19388,G19389,G19390,G19391,G19392,G19393,G19394,G19395,G19396,G19397,G19398,G19399,G19400,
       G19401,G19402,G19403,G19404,G19405,G19406,G19407,G19408,G19409,G19410,G19411,G19412,G19413,G19414,G19415,G19416,G19417,G19418,G19419,G19420,
       G19421,G19422,G19423,G19424,G19425,G19426,G19427,G19428,G19429,G19430,G19431,G19432,G19433,G19434,G19435,G19436,G19437,G19438,G19439,G19440,
       G19441,G19442,G19443,G19444,G19445,G19446,G19447,G19448,G19449,G19450,G19451,G19452,G19453,G19454,G19455,G19456,G19457,G19458,G19459,G19460,
       G19461,G19462,G19463,G19464,G19465,G19466,G19467,G19468,G19469,G19470,G19471,G19472,G19473,G19474,G19475,G19476,G19477,G19478,G19479,G19480,
       G19481,G19482,G19483,G19484,G19485,G19486,G19487,G19488,G19489,G19490,G19491,G19492,G19493,G19494,G19495,G19496,G19497,G19498,G19499,G19500,
       G19501,G19502,G19503,G19504,G19505,G19506,G19507,G19508,G19509,G19510,G19511,G19512,G19513,G19514,G19515,G19516,G19517,G19518,G19519,G19520,
       G19521,G19522,G19523,G19524,G19525,G19526,G19527,G19528,G19529,G19530,G19531,G19532,G19533,G19534,G19535,G19536,G19537,G19538,G19539,G19540,
       G19541,G19542,G19543,G19544,G19545,G19546,G19547,G19548,G19549,G19550,G19551,G19552,G19553,G19554,G19555,G19556,G19557,G19558,G19559,G19560,
       G19561,G19562,G19563,G19564,G19565,G19566,G19567,G19568,G19569,G19570,G19571,G19572,G19573,G19574,G19575,G19576,G19577,G19578,G19579,G19580,
       G19581,G19582,G19583,G19584,G19585,G19586,G19587,G19588,G19589,G19590,G19591,G19592,G19593,G19594,G19595,G19596,G19597,G19598,G19599,G19600,
       G19601,G19602,G19603,G19604,G19605,G19606,G19607,G19608,G19609,G19610,G19611,G19612,G19613,G19614,G19615,G19616,G19617,G19618,G19619,G19620,
       G19621,G19622,G19623,G19624,G19625,G19626,G19627,G19628,G19629,G19630,G19631,G19632,G19633,G19634,G19635,G19636,G19637,G19638,G19639,G19640,
       G19641,G19642,G19643,G19644,G19645,G19646,G19647,G19648,G19649,G19650,G19651,G19652,G19653,G19654,G19655,G19656,G19657,G19658,G19659,G19660,
       G19661,G19662,G19663,G19664,G19665,G19666,G19667,G19668,G19669,G19670,G19671,G19672,G19673,G19674,G19675,G19676,G19677,G19678,G19679,G19680,
       G19681,G19682,G19683,G19684,G19685,G19686,G19687,G19688,G19689,G19690,G19691,G19692,G19693,G19694,G19695,G19696,G19697,G19698,G19699,G19700,
       G19701,G19702,G19703,G19704,G19705,G19706,G19707,G19708,G19709,G19710,G19711,G19712,G19713,G19714,G19715,G19716,G19717,G19718,G19719,G19720,
       G19721,G19722,G19723,G19724,G19725,G19726,G19727,G19728,G19729,G19730,G19731,G19732,G19733,G19734,G19735,G19736,G19737,G19738,G19739,G19740,
       G19741,G19742,G19743,G19744,G19745,G19746,G19747,G19748,G19749,G19750,G19751,G19752,G19753,G19754,G19755,G19756,G19757,G19758,G19759,G19760,
       G19761,G19762,G19763,G19764,G19765,G19766,G19767,G19768,G19769,G19770,G19771,G19772,G19773,G19774,G19775,G19776,G19777,G19778,G19779,G19780,
       G19781,G19782,G19783,G19784,G19785,G19786,G19787,G19788,G19789,G19790,G19791,G19792,G19793,G19794,G19795,G19796,G19797,G19798,G19799,G19800,
       G19801,G19802,G19803,G19804,G19805,G19806,G19807,G19808,G19809,G19810,G19811,G19812,G19813,G19814,G19815,G19816,G19817,G19818,G19819,G19820,
       G19821,G19822,G19823,G19824,G19825,G19826,G19827,G19828,G19829,G19830,G19831,G19832,G19833,G19834,G19835,G19836,G19837,G19838,G19839,G19840,
       G19841,G19842,G19843,G19844,G19845,G19846,G19847,G19848,G19849,G19850,G19851,G19852,G19853,G19854,G19855,G19856,G19857,G19858,G19859,G19860,
       G19861,G19862,G19863,G19864,G19865,G19866,G19867,G19868,G19869,G19870,G19871,G19872,G19873,G19874,G19875,G19876,G19877,G19878,G19879,G19880,
       G19881,G19882,G19883,G19884,G19885,G19886,G19887,G19888,G19889,G19890,G19891,G19892,G19893,G19894,G19895,G19896,G19897,G19898,G19899,G19900,
       G19901,G19902,G19903,G19904,G19905,G19906,G19907,G19908,G19909,G19910,G19911,G19912,G19913,G19914,G19915,G19916,G19917,G19918,G19919,G19920,
       G19921,G19922,G19923,G19924,G19925,G19926,G19927,G19928,G19929,G19930,G19931,G19932,G19933,G19934,G19935,G19936,G19937,G19938,G19939,G19940,
       G19941,G19942,G19943,G19944,G19945,G19946,G19947,G19948,G19949,G19950,G19951,G19952,G19953,G19954,G19955,G19956,G19957,G19958,G19959,G19960,
       G19961,G19962,G19963,G19964,G19965,G19966,G19967,G19968,G19969,G19970,G19971,G19972,G19973,G19974,G19975,G19976,G19977,G19978,G19979,G19980,
       G19981,G19982,G19983,G19984,G19985,G19986,G19987,G19988,G19989,G19990,G19991,G19992,G19993,G19994,G19995,G19996,G19997,G19998,G19999,G20000,
       G20001,G20002,G20003,G20004,G20005,G20006,G20007,G20008,G20009,G20010,G20011,G20012,G20013,G20014,G20015,G20016,G20017,G20018,G20019,G20020,
       G20021,G20022,G20023,G20024,G20025,G20026,G20027,G20028,G20029,G20030,G20031,G20032,G20033,G20034,G20035,G20036,G20037,G20038,G20039,G20040,
       G20041,G20042,G20043,G20044,G20045,G20046,G20047,G20048,G20049,G20050,G20051,G20052,G20053,G20054,G20055,G20056,G20057,G20058,G20059,G20060,
       G20061,G20062,G20063,G20064,G20065,G20066,G20067,G20068,G20069,G20070,G20071,G20072,G20073,G20074,G20075,G20076,G20077,G20078,G20079,G20080,
       G20081,G20082,G20083,G20084,G20085,G20086,G20087,G20088,G20089,G20090,G20091,G20092,G20093,G20094,G20095,G20096,G20097,G20098,G20099,G20100,
       G20101,G20102,G20103,G20104,G20105,G20106,G20107,G20108,G20109,G20110,G20111,G20112,G20113,G20114,G20115,G20116,G20117,G20118,G20119,G20120,
       G20121,G20122,G20123,G20124,G20125,G20126,G20127,G20128,G20129,G20130,G20131,G20132,G20133,G20134,G20135,G20136,G20137,G20138,G20139,G20140,
       G20141,G20142,G20143,G20144,G20145,G20146,G20147,G20148,G20149,G20150,G20151,G20152,G20153,G20154,G20155,G20156,G20157,G20158,G20159,G20160,
       G20161,G20162,G20163,G20164,G20165,G20166,G20167,G20168,G20169,G20170,G20171,G20172,G20173,G20174,G20175,G20176,G20177,G20178,G20179,G20180,
       G20181,G20182,G20183,G20184,G20185,G20186,G20187,G20188,G20189,G20190,G20191,G20192,G20193,G20194,G20195,G20196,G20197,G20198,G20199,G20200,
       G20201,G20202,G20203,G20204,G20205,G20206,G20207,G20208,G20209,G20210,G20211,G20212,G20213,G20214,G20215,G20216,G20217,G20218,G20219,G20220,
       G20221,G20222,G20223,G20224,G20225,G20226,G20227,G20228,G20229,G20230,G20231,G20232,G20233,G20234,G20235,G20236,G20237,G20238,G20239,G20240,
       G20241,G20242,G20243,G20244,G20245,G20246,G20247,G20248,G20249,G20250,G20251,G20252,G20253,G20254,G20255,G20256,G20257,G20258,G20259,G20260,
       G20261,G20262,G20263,G20264,G20265,G20266,G20267,G20268,G20269,G20270,G20271,G20272,G20273,G20274,G20275,G20276,G20277,G20278,G20279,G20280,
       G20281,G20282,G20283,G20284,G20285,G20286,G20287,G20288,G20289,G20290,G20291,G20292,G20293,G20294,G20295,G20296,G20297,G20298,G20299,G20300,
       G20301,G20302,G20303,G20304,G20305,G20306,G20307,G20308,G20309,G20310,G20311,G20312,G20313,G20314,G20315,G20316,G20317,G20318,G20319,G20320,
       G20321,G20322,G20323,G20324,G20325,G20326,G20327,G20328,G20329,G20330,G20331,G20332,G20333,G20334,G20335,G20336,G20337,G20338,G20339,G20340,
       G20341,G20342,G20343,G20344,G20345,G20346,G20347,G20348,G20349,G20350,G20351,G20352,G20353,G20354,G20355,G20356,G20357,G20358,G20359,G20360,
       G20361,G20362,G20363,G20364,G20365,G20366,G20367,G20368,G20369,G20370,G20371,G20372,G20373,G20374,G20375,G20376,G20377,G20378,G20379,G20380,
       G20381,G20382,G20383,G20384,G20385,G20386,G20387,G20388,G20389,G20390,G20391,G20392,G20393,G20394,G20395,G20396,G20397,G20398,G20399,G20400,
       G20401,G20402,G20403,G20404,G20405,G20406,G20407,G20408,G20409,G20410,G20411,G20412,G20413,G20414,G20415,G20416,G20417,G20418,G20419,G20420,
       G20421,G20422,G20423,G20424,G20425,G20426,G20427,G20428,G20429,G20430,G20431,G20432,G20433,G20434,G20435,G20436,G20437,G20438,G20439,G20440,
       G20441,G20442,G20443,G20444,G20445,G20446,G20447,G20448,G20449,G20450,G20451,G20452,G20453,G20454,G20455,G20456,G20457,G20458,G20459,G20460,
       G20461,G20462,G20463,G20464,G20465,G20466,G20467,G20468,G20469,G20470,G20471,G20472,G20473,G20474,G20475,G20476,G20477,G20478,G20479,G20480,
       G20481,G20482,G20483,G20484,G20485,G20486,G20487,G20488,G20489,G20490,G20491,G20492,G20493,G20494,G20495,G20496,G20497,G20498,G20499,G20500,
       G20501,G20502,G20503,G20504,G20505,G20506,G20507,G20508,G20509,G20510,G20511,G20512,G20513,G20514,G20515,G20516,G20517,G20518,G20519,G20520,
       G20521,G20522,G20523,G20524,G20525,G20526,G20527,G20528,G20529,G20530,G20531,G20532,G20533,G20534,G20535,G20536,G20537,G20538,G20539,G20540,
       G20541,G20542,G20543,G20544,G20545,G20546,G20547,G20548,G20549,G20550,G20551,G20552,G20553,G20554,G20555,G20556,G20557,G20558,G20559,G20560,
       G20561,G20562,G20563,G20564,G20565,G20566,G20567,G20568,G20569,G20570,G20571,G20572,G20573,G20574,G20575,G20576,G20577,G20578,G20579,G20580,
       G20581,G20582,G20583,G20584,G20585,G20586,G20587,G20588,G20589,G20590,G20591,G20592,G20593,G20594,G20595,G20596,G20597,G20598,G20599,G20600,
       G20601,G20602,G20603,G20604,G20605,G20606,G20607,G20608,G20609,G20610,G20611,G20612,G20613,G20614,G20615,G20616,G20617,G20618,G20619,G20620,
       G20621,G20622,G20623,G20624,G20625,G20626,G20627,G20628,G20629,G20630,G20631,G20632,G20633,G20634,G20635,G20636,G20637,G20638,G20639,G20640,
       G20641,G20642,G20643,G20644,G20645,G20646,G20647,G20648,G20649,G20650,G20651,G20652,G20653,G20654,G20655,G20656,G20657,G20658,G20659,G20660,
       G20661,G20662,G20663,G20664,G20665,G20666,G20667,G20668,G20669,G20670,G20671,G20672,G20673,G20674,G20675,G20676,G20677,G20678,G20679,G20680,
       G20681,G20682,G20683,G20684,G20685,G20686,G20687,G20688,G20689,G20690,G20691,G20692,G20693,G20694,G20695,G20696,G20697,G20698,G20699,G20700,
       G20701,G20702,G20703,G20704,G20705,G20706,G20707,G20708,G20709,G20710,G20711,G20712,G20713,G20714,G20715,G20716,G20717,G20718,G20719,G20720,
       G20721,G20722,G20723,G20724,G20725,G20726,G20727,G20728,G20729,G20730,G20731,G20732,G20733,G20734,G20735,G20736,G20737,G20738,G20739,G20740,
       G20741,G20742,G20743,G20744,G20745,G20746,G20747,G20748,G20749,G20750,G20751,G20752,G20753,G20754,G20755,G20756,G20757,G20758,G20759,G20760,
       G20761,G20762,G20763,G20764,G20765,G20766,G20767,G20768,G20769,G20770,G20771,G20772,G20773,G20774,G20775,G20776,G20777,G20778,G20779,G20780,
       G20781,G20782,G20783,G20784,G20785,G20786,G20787,G20788,G20789,G20790,G20791,G20792,G20793,G20794,G20795,G20796,G20797,G20798,G20799,G20800,
       G20801,G20802,G20803,G20804,G20805,G20806,G20807,G20808,G20809,G20810,G20811,G20812,G20813,G20814,G20815,G20816,G20817,G20818,G20819,G20820,
       G20821,G20822,G20823,G20824,G20825,G20826,G20827,G20828,G20829,G20830,G20831,G20832,G20833,G20834,G20835,G20836,G20837,G20838,G20839,G20840,
       G20841,G20842,G20843,G20844,G20845,G20846,G20847,G20848,G20849,G20850,G20851,G20852,G20853,G20854,G20855,G20856,G20857,G20858,G20859,G20860,
       G20861,G20862,G20863,G20864,G20865,G20866,G20867,G20868,G20869,G20870,G20871,G20872,G20873,G20874,G20875,G20876,G20877,G20878,G20879,G20880,
       G20881,G20882,G20883,G20884,G20885,G20886,G20887,G20888,G20889,G20890,G20891,G20892,G20893,G20894,G20895,G20896,G20897,G20898,G20899,G20900,
       G20901,G20902,G20903,G20904,G20905,G20906,G20907,G20908,G20909,G20910,G20911,G20912,G20913,G20914,G20915,G20916,G20917,G20918,G20919,G20920,
       G20921,G20922,G20923,G20924,G20925,G20926,G20927,G20928,G20929,G20930,G20931,G20932,G20933,G20934,G20935,G20936,G20937,G20938,G20939,G20940,
       G20941,G20942,G20943,G20944,G20945,G20946,G20947,G20948,G20949,G20950,G20951,G20952,G20953,G20954,G20955,G20956,G20957,G20958,G20959,G20960,
       G20961,G20962,G20963,G20964,G20965,G20966,G20967,G20968,G20969,G20970,G20971,G20972,G20973,G20974,G20975,G20976,G20977,G20978,G20979,G20980,
       G20981,G20982,G20983,G20984,G20985,G20986,G20987,G20988,G20989,G20990,G20991,G20992,G20993,G20994,G20995,G20996,G20997,G20998,G20999,G21000,
       G21001,G21002,G21003,G21004,G21005,G21006,G21007,G21008,G21009,G21010,G21011,G21012,G21013,G21014,G21015,G21016,G21017,G21018,G21019,G21020,
       G21021,G21022,G21023,G21024,G21025,G21026,G21027,G21028,G21029,G21030,G21031,G21032,G21033,G21034,G21035,G21036,G21037,G21038,G21039,G21040,
       G21041,G21042,G21043,G21044,G21045,G21046,G21047,G21048,G21049,G21050,G21051,G21052,G21053,G21054,G21055,G21056,G21057,G21058,G21059,G21060,
       G21061,G21062,G21063,G21064,G21065,G21066,G21067,G21068,G21069,G21070,G21071,G21072,G21073,G21074,G21075,G21076,G21077,G21078,G21079,G21080,
       G21081,G21082,G21083,G21084,G21085,G21086,G21087,G21088,G21089,G21090,G21091,G21092,G21093,G21094,G21095,G21096,G21097,G21098,G21099,G21100,
       G21101,G21102,G21103,G21104,G21105,G21106,G21107,G21108,G21109,G21110,G21111,G21112,G21113,G21114,G21115,G21116,G21117,G21118,G21119,G21120,
       G21121,G21122,G21123,G21124,G21125,G21126,G21127,G21128,G21129,G21130,G21131,G21132,G21133,G21134,G21135,G21136,G21137,G21138,G21139,G21140,
       G21141,G21142,G21143,G21144,G21145,G21146,G21147,G21148,G21149,G21150,G21151,G21152,G21153,G21154,G21155,G21156,G21157,G21158,G21159,G21160,
       G21161,G21162,G21163,G21164,G21165,G21166,G21167,G21168,G21169,G21170,G21171,G21172,G21173,G21174,G21175,G21176,G21177,G21178,G21179,G21180,
       G21181,G21182,G21183,G21184,G21185,G21186,G21187,G21188,G21189,G21190,G21191,G21192,G21193,G21194,G21195,G21196,G21197,G21198,G21199,G21200,
       G21201,G21202,G21203,G21204,G21205,G21206,G21207,G21208,G21209,G21210,G21211,G21212,G21213,G21214,G21215,G21216,G21217,G21218,G21219,G21220,
       G21221,G21222,G21223,G21224,G21225,G21226,G21227,G21228,G21229,G21230,G21231,G21232,G21233,G21234,G21235,G21236,G21237,G21238,G21239,G21240,
       G21241,G21242,G21243,G21244,G21245,G21246,G21247,G21248,G21249,G21250,G21251,G21252,G21253,G21254,G21255,G21256,G21257,G21258,G21259,G21260,
       G21261,G21262,G21263,G21264,G21265,G21266,G21267,G21268,G21269,G21270,G21271,G21272,G21273,G21274,G21275,G21276,G21277,G21278,G21279,G21280,
       G21281,G21282,G21283,G21284,G21285,G21286,G21287,G21288,G21289,G21290,G21291,G21292,G21293,G21294,G21295,G21296,G21297,G21298,G21299,G21300,
       G21301,G21302,G21303,G21304,G21305,G21306,G21307,G21308,G21309,G21310,G21311,G21312,G21313,G21314,G21315,G21316,G21317,G21318,G21319,G21320,
       G21321,G21322,G21323,G21324,G21325,G21326,G21327,G21328,G21329,G21330,G21331,G21332,G21333,G21334,G21335,G21336,G21337,G21338,G21339,G21340,
       G21341,G21342,G21343,G21344,G21345,G21346,G21347,G21348,G21349,G21350,G21351,G21352,G21353,G21354,G21355,G21356,G21357,G21358,G21359,G21360,
       G21361,G21362,G21363,G21364,G21365,G21366,G21367,G21368,G21369,G21370,G21371,G21372,G21373,G21374,G21375,G21376,G21377,G21378,G21379,G21380,
       G21381,G21382,G21383,G21384,G21385,G21386,G21387,G21388,G21389,G21390,G21391,G21392,G21393,G21394,G21395,G21396,G21397,G21398,G21399,G21400,
       G21401,G21402,G21403,G21404,G21405,G21406,G21407,G21408,G21409,G21410,G21411,G21412,G21413,G21414,G21415,G21416,G21417,G21418,G21419,G21420,
       G21421,G21422,G21423,G21424,G21425,G21426,G21427,G21428,G21429,G21430,G21431,G21432,G21433,G21434,G21435,G21436,G21437,G21438,G21439,G21440,
       G21441,G21442,G21443,G21444,G21445,G21446,G21447,G21448,G21449,G21450,G21451,G21452,G21453,G21454,G21455,G21456,G21457,G21458,G21459,G21460,
       G21461,G21462,G21463,G21464,G21465,G21466,G21467,G21468,G21469,G21470,G21471,G21472,G21473,G21474,G21475,G21476,G21477,G21478,G21479,G21480,
       G21481,G21482,G21483,G21484,G21485,G21486,G21487,G21488,G21489,G21490,G21491,G21492,G21493,G21494,G21495,G21496,G21497,G21498,G21499,G21500,
       G21501,G21502,G21503,G21504,G21505,G21506,G21507,G21508,G21509,G21510,G21511,G21512,G21513,G21514,G21515,G21516,G21517,G21518,G21519,G21520,
       G21521,G21522,G21523,G21524,G21525,G21526,G21527,G21528,G21529,G21530,G21531,G21532,G21533,G21534,G21535,G21536,G21537,G21538,G21539,G21540,
       G21541,G21542,G21543,G21544,G21545,G21546,G21547,G21548,G21549,G21550,G21551,G21552,G21553,G21554,G21555,G21556,G21557,G21558,G21559,G21560,
       G21561,G21562,G21563,G21564,G21565,G21566,G21567,G21568,G21569,G21570,G21571,G21572,G21573,G21574,G21575,G21576,G21577,G21578,G21579,G21580,
       G21581,G21582,G21583,G21584,G21585,G21586,G21587,G21588,G21589,G21590,G21591,G21592,G21593,G21594,G21595,G21596,G21597,G21598,G21599,G21600,
       G21601,G21602,G21603,G21604,G21605,G21606,G21607,G21608,G21609,G21610,G21611,G21612,G21613,G21614,G21615,G21616,G21617,G21618,G21619,G21620,
       G21621,G21622,G21623,G21624,G21625,G21626,G21627,G21628,G21629,G21630,G21631,G21632,G21633,G21634,G21635,G21636,G21637,G21638,G21639,G21640,
       G21641,G21642,G21643,G21644,G21645,G21646,G21647,G21648,G21649,G21650,G21651,G21652,G21653,G21654,G21655,G21656,G21657,G21658,G21659,G21660,
       G21661,G21662,G21663,G21664,G21665,G21666,G21667,G21668,G21669,G21670,G21671,G21672,G21673,G21674,G21675,G21676,G21677,G21678,G21679,G21680,
       G21681,G21682,G21683,G21684,G21685,G21686,G21687,G21688,G21689,G21690,G21691,G21692,G21693,G21694,G21695,G21696,G21697,G21698,G21699,G21700,
       G21701,G21702,G21703,G21704,G21705,G21706,G21707,G21708,G21709,G21710,G21711,G21712,G21713,G21714,G21715,G21716,G21717,G21718,G21719,G21720,
       G21721,G21722,G21723,G21724,G21725,G21726,G21727,G21728,G21729,G21730,G21731,G21732,G21733,G21734,G21735,G21736,G21737,G21738,G21739,G21740,
       G21741,G21742,G21743,G21744,G21745,G21746,G21747,G21748,G21749,G21750,G21751,G21752,G21753,G21754,G21755,G21756,G21757,G21758,G21759,G21760,
       G21761,G21762,G21763,G21764,G21765,G21766,G21767,G21768,G21769,G21770,G21771,G21772,G21773,G21774,G21775,G21776,G21777,G21778,G21779,G21780,
       G21781,G21782,G21783,G21784,G21785,G21786,G21787,G21788,G21789,G21790,G21791,G21792,G21793,G21794,G21795,G21796,G21797,G21798,G21799,G21800,
       G21801,G21802,G21803,G21804;

  dff DFF_107(CK,G21356,G1732);
  dff DFF_108(CK,G21357,G1733);
  dff DFF_109(CK,G21358,G1734);
  dff DFF_110(CK,G21359,G1735);
  dff DFF_111(CK,G21360,G757);
  dff DFF_112(CK,G21361,G758);
  dff DFF_113(CK,G21362,G759);
  dff DFF_114(CK,G21363,G760);
  dff DFF_115(CK,G21364,G761);
  dff DFF_116(CK,G21365,G762);
  dff DFF_117(CK,G21366,G763);
  dff DFF_118(CK,G21367,G764);
  dff DFF_119(CK,G21368,G765);
  dff DFF_120(CK,G21369,G766);
  dff DFF_121(CK,G21370,G767);
  dff DFF_122(CK,G21371,G768);
  dff DFF_123(CK,G21372,G769);
  dff DFF_124(CK,G21373,G770);
  dff DFF_125(CK,G21374,G771);
  dff DFF_126(CK,G21375,G772);
  dff DFF_127(CK,G21376,G773);
  dff DFF_128(CK,G21377,G774);
  dff DFF_129(CK,G21378,G775);
  dff DFF_130(CK,G21379,G776);
  dff DFF_131(CK,G21380,G777);
  dff DFF_132(CK,G21381,G778);
  dff DFF_133(CK,G21382,G779);
  dff DFF_134(CK,G21383,G780);
  dff DFF_135(CK,G21384,G781);
  dff DFF_136(CK,G21385,G782);
  dff DFF_137(CK,G21386,G783);
  dff DFF_138(CK,G21387,G784);
  dff DFF_139(CK,G21388,G785);
  dff DFF_140(CK,G21389,G786);
  dff DFF_141(CK,G21390,G787);
  dff DFF_142(CK,G21391,G789);
  dff DFF_143(CK,G21392,G790);
  dff DFF_144(CK,G21393,G1737);
  dff DFF_145(CK,G21394,G1738);
  dff DFF_146(CK,G21395,G791);
  dff DFF_147(CK,G21396,G792);
  dff DFF_148(CK,G21397,G793);
  dff DFF_149(CK,G21398,G794);
  dff DFF_150(CK,G21399,G795);
  dff DFF_151(CK,G21400,G796);
  dff DFF_152(CK,G21401,G797);
  dff DFF_153(CK,G21402,G798);
  dff DFF_154(CK,G21403,G799);
  dff DFF_155(CK,G21404,G800);
  dff DFF_156(CK,G21405,G801);
  dff DFF_157(CK,G21406,G802);
  dff DFF_158(CK,G21407,G803);
  dff DFF_159(CK,G21408,G804);
  dff DFF_160(CK,G21409,G805);
  dff DFF_161(CK,G21410,G806);
  dff DFF_162(CK,G21411,G807);
  dff DFF_163(CK,G21412,G808);
  dff DFF_164(CK,G21413,G809);
  dff DFF_165(CK,G21414,G810);
  dff DFF_166(CK,G21415,G811);
  dff DFF_167(CK,G21416,G812);
  dff DFF_168(CK,G21417,G813);
  dff DFF_169(CK,G21418,G814);
  dff DFF_170(CK,G21419,G815);
  dff DFF_171(CK,G21420,G816);
  dff DFF_172(CK,G21421,G817);
  dff DFF_173(CK,G21422,G818);
  dff DFF_174(CK,G21423,G819);
  dff DFF_175(CK,G21424,G820);
  dff DFF_176(CK,G21425,G821);
  dff DFF_177(CK,G21426,G822);
  dff DFF_178(CK,G21427,G823);
  dff DFF_179(CK,G21428,G824);
  dff DFF_180(CK,G21429,G825);
  dff DFF_181(CK,G21430,G826);
  dff DFF_182(CK,G21431,G827);
  dff DFF_183(CK,G21432,G828);
  dff DFF_184(CK,G21433,G829);
  dff DFF_185(CK,G21434,G830);
  dff DFF_186(CK,G21435,G831);
  dff DFF_187(CK,G21436,G832);
  dff DFF_188(CK,G21437,G833);
  dff DFF_189(CK,G21438,G834);
  dff DFF_190(CK,G21439,G835);
  dff DFF_191(CK,G21440,G836);
  dff DFF_192(CK,G21441,G837);
  dff DFF_193(CK,G21442,G838);
  dff DFF_194(CK,G21443,G839);
  dff DFF_195(CK,G21444,G840);
  dff DFF_196(CK,G21445,G841);
  dff DFF_197(CK,G21446,G842);
  dff DFF_198(CK,G21447,G843);
  dff DFF_199(CK,G21448,G844);
  dff DFF_200(CK,G21449,G845);
  dff DFF_201(CK,G21450,G846);
  dff DFF_202(CK,G21451,G847);
  dff DFF_203(CK,G21452,G848);
  dff DFF_204(CK,G21453,G849);
  dff DFF_205(CK,G21454,G850);
  dff DFF_206(CK,G21455,G851);
  dff DFF_207(CK,G21456,G852);
  dff DFF_208(CK,G21457,G853);
  dff DFF_209(CK,G21458,G854);
  dff DFF_210(CK,G21459,G855);
  dff DFF_211(CK,G21460,G856);
  dff DFF_212(CK,G21461,G857);
  dff DFF_213(CK,G21462,G858);
  dff DFF_214(CK,G21463,G859);
  dff DFF_215(CK,G21464,G860);
  dff DFF_216(CK,G21465,G861);
  dff DFF_217(CK,G21466,G862);
  dff DFF_218(CK,G21467,G863);
  dff DFF_219(CK,G21468,G864);
  dff DFF_220(CK,G21469,G865);
  dff DFF_221(CK,G21470,G866);
  dff DFF_222(CK,G21471,G867);
  dff DFF_223(CK,G21472,G868);
  dff DFF_224(CK,G21473,G869);
  dff DFF_225(CK,G21474,G870);
  dff DFF_226(CK,G21475,G871);
  dff DFF_227(CK,G21476,G872);
  dff DFF_228(CK,G21477,G873);
  dff DFF_229(CK,G21478,G874);
  dff DFF_230(CK,G21479,G875);
  dff DFF_231(CK,G21480,G876);
  dff DFF_232(CK,G21481,G877);
  dff DFF_233(CK,G21482,G878);
  dff DFF_234(CK,G21483,G879);
  dff DFF_235(CK,G21484,G880);
  dff DFF_236(CK,G21485,G881);
  dff DFF_237(CK,G21486,G882);
  dff DFF_238(CK,G21487,G883);
  dff DFF_239(CK,G21488,G884);
  dff DFF_240(CK,G21489,G885);
  dff DFF_241(CK,G21490,G886);
  dff DFF_242(CK,G21491,G887);
  dff DFF_243(CK,G21492,G888);
  dff DFF_244(CK,G21493,G889);
  dff DFF_245(CK,G21494,G890);
  dff DFF_246(CK,G21495,G891);
  dff DFF_247(CK,G21496,G892);
  dff DFF_248(CK,G21497,G893);
  dff DFF_249(CK,G21498,G894);
  dff DFF_250(CK,G21499,G895);
  dff DFF_251(CK,G21500,G896);
  dff DFF_252(CK,G21501,G897);
  dff DFF_253(CK,G21502,G898);
  dff DFF_254(CK,G21503,G899);
  dff DFF_255(CK,G21504,G900);
  dff DFF_256(CK,G21505,G901);
  dff DFF_257(CK,G21506,G902);
  dff DFF_258(CK,G21507,G903);
  dff DFF_259(CK,G21508,G904);
  dff DFF_260(CK,G21509,G905);
  dff DFF_261(CK,G21510,G906);
  dff DFF_262(CK,G21511,G907);
  dff DFF_263(CK,G21512,G908);
  dff DFF_264(CK,G21513,G909);
  dff DFF_265(CK,G21514,G910);
  dff DFF_266(CK,G21515,G911);
  dff DFF_267(CK,G21516,G912);
  dff DFF_268(CK,G21517,G913);
  dff DFF_269(CK,G21518,G914);
  dff DFF_270(CK,G21519,G915);
  dff DFF_271(CK,G21520,G916);
  dff DFF_272(CK,G21521,G917);
  dff DFF_273(CK,G21522,G918);
  dff DFF_274(CK,G21523,G919);
  dff DFF_275(CK,G21524,G920);
  dff DFF_276(CK,G21525,G921);
  dff DFF_277(CK,G21526,G922);
  dff DFF_278(CK,G21527,G923);
  dff DFF_279(CK,G21528,G924);
  dff DFF_280(CK,G21529,G925);
  dff DFF_281(CK,G21530,G926);
  dff DFF_282(CK,G21531,G927);
  dff DFF_283(CK,G21532,G928);
  dff DFF_284(CK,G21533,G929);
  dff DFF_285(CK,G21534,G930);
  dff DFF_286(CK,G21535,G931);
  dff DFF_287(CK,G21536,G932);
  dff DFF_288(CK,G21537,G933);
  dff DFF_289(CK,G21538,G934);
  dff DFF_290(CK,G21539,G935);
  dff DFF_291(CK,G21540,G936);
  dff DFF_292(CK,G21541,G937);
  dff DFF_293(CK,G21542,G938);
  dff DFF_294(CK,G21543,G939);
  dff DFF_295(CK,G21544,G940);
  dff DFF_296(CK,G21545,G941);
  dff DFF_297(CK,G21546,G942);
  dff DFF_298(CK,G21547,G943);
  dff DFF_299(CK,G21548,G944);
  dff DFF_300(CK,G21549,G945);
  dff DFF_301(CK,G21550,G946);
  dff DFF_302(CK,G21551,G947);
  dff DFF_303(CK,G21552,G948);
  dff DFF_304(CK,G21553,G949);
  dff DFF_305(CK,G21554,G950);
  dff DFF_306(CK,G21555,G951);
  dff DFF_307(CK,G21556,G952);
  dff DFF_308(CK,G21557,G1740);
  dff DFF_309(CK,G21558,G1742);
  dff DFF_310(CK,G21559,G1743);
  dff DFF_311(CK,G21560,G1744);
  dff DFF_312(CK,G21561,G1745);
  dff DFF_313(CK,G21562,G953);
  dff DFF_314(CK,G21563,G954);
  dff DFF_315(CK,G21564,G955);
  dff DFF_316(CK,G21565,G956);
  dff DFF_317(CK,G21566,G1746);
  dff DFF_318(CK,G21567,G957);
  dff DFF_319(CK,G21568,G958);
  dff DFF_320(CK,G21569,G959);
  dff DFF_321(CK,G21570,G960);
  dff DFF_322(CK,G21571,G961);
  dff DFF_323(CK,G21572,G962);
  dff DFF_324(CK,G21573,G963);
  dff DFF_325(CK,G21574,G964);
  dff DFF_326(CK,G21575,G965);
  dff DFF_327(CK,G21576,G966);
  dff DFF_328(CK,G21577,G967);
  dff DFF_329(CK,G21578,G968);
  dff DFF_330(CK,G21579,G969);
  dff DFF_331(CK,G21580,G970);
  dff DFF_332(CK,G21581,G971);
  dff DFF_333(CK,G21582,G972);
  dff DFF_334(CK,G21583,G973);
  dff DFF_335(CK,G21584,G974);
  dff DFF_336(CK,G21585,G975);
  dff DFF_337(CK,G21586,G976);
  dff DFF_338(CK,G21587,G977);
  dff DFF_339(CK,G21588,G978);
  dff DFF_340(CK,G21589,G979);
  dff DFF_341(CK,G21590,G980);
  dff DFF_342(CK,G21591,G981);
  dff DFF_343(CK,G21592,G982);
  dff DFF_344(CK,G21593,G983);
  dff DFF_345(CK,G21594,G984);
  dff DFF_346(CK,G21595,G985);
  dff DFF_347(CK,G21596,G986);
  dff DFF_348(CK,G21597,G987);
  dff DFF_349(CK,G21598,G988);
  dff DFF_350(CK,G21599,G989);
  dff DFF_351(CK,G21600,G990);
  dff DFF_352(CK,G21601,G991);
  dff DFF_353(CK,G21602,G992);
  dff DFF_354(CK,G21603,G993);
  dff DFF_355(CK,G21604,G994);
  dff DFF_356(CK,G21605,G995);
  dff DFF_357(CK,G21606,G996);
  dff DFF_358(CK,G21607,G997);
  dff DFF_359(CK,G21608,G998);
  dff DFF_360(CK,G21609,G999);
  dff DFF_361(CK,G21610,G1000);
  dff DFF_362(CK,G21611,G1001);
  dff DFF_363(CK,G21612,G1002);
  dff DFF_364(CK,G21613,G1003);
  dff DFF_365(CK,G21614,G1004);
  dff DFF_366(CK,G21615,G1005);
  dff DFF_367(CK,G21616,G1006);
  dff DFF_368(CK,G21617,G1007);
  dff DFF_369(CK,G21618,G1008);
  dff DFF_370(CK,G21619,G1009);
  dff DFF_371(CK,G21620,G1010);
  dff DFF_372(CK,G21621,G1011);
  dff DFF_373(CK,G21622,G1012);
  dff DFF_374(CK,G21623,G1013);
  dff DFF_375(CK,G21624,G1014);
  dff DFF_376(CK,G21625,G1015);
  dff DFF_377(CK,G21626,G1016);
  dff DFF_378(CK,G21627,G1017);
  dff DFF_379(CK,G21628,G1018);
  dff DFF_380(CK,G21629,G1019);
  dff DFF_381(CK,G21630,G1020);
  dff DFF_382(CK,G21631,G1021);
  dff DFF_383(CK,G21632,G1022);
  dff DFF_384(CK,G21633,G1023);
  dff DFF_385(CK,G21634,G1024);
  dff DFF_386(CK,G21635,G1025);
  dff DFF_387(CK,G21636,G1026);
  dff DFF_388(CK,G21637,G1027);
  dff DFF_389(CK,G21638,G1028);
  dff DFF_390(CK,G21639,G1029);
  dff DFF_391(CK,G21640,G1030);
  dff DFF_392(CK,G21641,G1031);
  dff DFF_393(CK,G21642,G1032);
  dff DFF_394(CK,G21643,G1033);
  dff DFF_395(CK,G21644,G1034);
  dff DFF_396(CK,G21645,G1035);
  dff DFF_397(CK,G21646,G1036);
  dff DFF_398(CK,G21647,G1037);
  dff DFF_399(CK,G21648,G1038);
  dff DFF_400(CK,G21649,G1039);
  dff DFF_401(CK,G21650,G1040);
  dff DFF_402(CK,G21651,G1041);
  dff DFF_403(CK,G21652,G1042);
  dff DFF_404(CK,G21653,G1043);
  dff DFF_405(CK,G21654,G1044);
  dff DFF_406(CK,G21655,G1045);
  dff DFF_407(CK,G21656,G1046);
  dff DFF_408(CK,G21657,G1047);
  dff DFF_409(CK,G21658,G1048);
  dff DFF_410(CK,G21659,G1049);
  dff DFF_411(CK,G21660,G1050);
  dff DFF_412(CK,G21661,G1051);
  dff DFF_413(CK,G21662,G1052);
  dff DFF_414(CK,G21663,G1053);
  dff DFF_415(CK,G21664,G1054);
  dff DFF_416(CK,G21665,G1055);
  dff DFF_417(CK,G21666,G1056);
  dff DFF_418(CK,G21667,G1057);
  dff DFF_419(CK,G21668,G1058);
  dff DFF_420(CK,G21669,G1059);
  dff DFF_421(CK,G21670,G1060);
  dff DFF_422(CK,G21671,G1061);
  dff DFF_423(CK,G21672,G1062);
  dff DFF_424(CK,G21673,G1063);
  dff DFF_425(CK,G21674,G1064);
  dff DFF_426(CK,G21675,G1065);
  dff DFF_427(CK,G21676,G1066);
  dff DFF_428(CK,G21677,G1067);
  dff DFF_429(CK,G21678,G1068);
  dff DFF_430(CK,G21679,G1069);
  dff DFF_431(CK,G21680,G1070);
  dff DFF_432(CK,G21681,G1071);
  dff DFF_433(CK,G21682,G1072);
  dff DFF_434(CK,G21683,G1073);
  dff DFF_435(CK,G21684,G1074);
  dff DFF_436(CK,G21685,G1075);
  dff DFF_437(CK,G21686,G1076);
  dff DFF_438(CK,G21687,G1077);
  dff DFF_439(CK,G21688,G1078);
  dff DFF_440(CK,G21689,G1079);
  dff DFF_441(CK,G21690,G1080);
  dff DFF_442(CK,G21691,G1081);
  dff DFF_443(CK,G21692,G1082);
  dff DFF_444(CK,G21693,G1083);
  dff DFF_445(CK,G21694,G1084);
  dff DFF_446(CK,G21695,G1085);
  dff DFF_447(CK,G21696,G1086);
  dff DFF_448(CK,G21697,G1087);
  dff DFF_449(CK,G21698,G1088);
  dff DFF_450(CK,G21699,G1089);
  dff DFF_451(CK,G21700,G1090);
  dff DFF_452(CK,G21701,G1091);
  dff DFF_453(CK,G21702,G1092);
  dff DFF_454(CK,G21703,G1093);
  dff DFF_455(CK,G21704,G1094);
  dff DFF_456(CK,G21705,G1095);
  dff DFF_457(CK,G21706,G1096);
  dff DFF_458(CK,G21707,G1097);
  dff DFF_459(CK,G21708,G1098);
  dff DFF_460(CK,G21709,G1099);
  dff DFF_461(CK,G21710,G1100);
  dff DFF_462(CK,G21711,G1101);
  dff DFF_463(CK,G21712,G1102);
  dff DFF_464(CK,G21713,G1103);
  dff DFF_465(CK,G21714,G1104);
  dff DFF_466(CK,G21715,G1105);
  dff DFF_467(CK,G21716,G1106);
  dff DFF_468(CK,G21717,G1107);
  dff DFF_469(CK,G21718,G1108);
  dff DFF_470(CK,G21719,G1109);
  dff DFF_471(CK,G21720,G1110);
  dff DFF_472(CK,G21721,G1111);
  dff DFF_473(CK,G21722,G1112);
  dff DFF_474(CK,G21723,G1113);
  dff DFF_475(CK,G21724,G1114);
  dff DFF_476(CK,G21725,G1115);
  dff DFF_477(CK,G21726,G1116);
  dff DFF_478(CK,G21727,G1117);
  dff DFF_479(CK,G21728,G1118);
  dff DFF_480(CK,G21729,G1119);
  dff DFF_481(CK,G21730,G1120);
  dff DFF_482(CK,G21731,G1121);
  dff DFF_483(CK,G21732,G1122);
  dff DFF_484(CK,G21733,G1123);
  dff DFF_485(CK,G21734,G1124);
  dff DFF_486(CK,G21735,G1125);
  dff DFF_487(CK,G21736,G1126);
  dff DFF_488(CK,G21737,G1127);
  dff DFF_489(CK,G21738,G1128);
  dff DFF_490(CK,G21739,G1129);
  dff DFF_491(CK,G21740,G1130);
  dff DFF_492(CK,G21741,G1131);
  dff DFF_493(CK,G21742,G1132);
  dff DFF_494(CK,G21743,G1133);
  dff DFF_495(CK,G21744,G1134);
  dff DFF_496(CK,G21745,G1135);
  dff DFF_497(CK,G21746,G1136);
  dff DFF_498(CK,G21747,G1137);
  dff DFF_499(CK,G21748,G1138);
  dff DFF_500(CK,G21749,G1139);
  dff DFF_501(CK,G21750,G1140);
  dff DFF_502(CK,G21751,G1141);
  dff DFF_503(CK,G21752,G1142);
  dff DFF_504(CK,G21753,G1143);
  dff DFF_505(CK,G21754,G1144);
  dff DFF_506(CK,G21755,G1145);
  dff DFF_507(CK,G21756,G1146);
  dff DFF_508(CK,G21757,G1147);
  dff DFF_509(CK,G21758,G1148);
  dff DFF_510(CK,G21759,G1149);
  dff DFF_511(CK,G21760,G1150);
  dff DFF_512(CK,G21761,G1151);
  dff DFF_513(CK,G21762,G1152);
  dff DFF_514(CK,G21763,G1153);
  dff DFF_515(CK,G21764,G1154);
  dff DFF_516(CK,G21765,G1155);
  dff DFF_517(CK,G21766,G1156);
  dff DFF_518(CK,G21767,G1157);
  dff DFF_519(CK,G21768,G1158);
  dff DFF_520(CK,G21769,G1159);
  dff DFF_521(CK,G21770,G1160);
  dff DFF_522(CK,G21771,G1161);
  dff DFF_523(CK,G21772,G1162);
  dff DFF_524(CK,G21773,G1163);
  dff DFF_525(CK,G21774,G1164);
  dff DFF_526(CK,G21775,G1165);
  dff DFF_527(CK,G21776,G1166);
  dff DFF_528(CK,G21777,G1167);
  dff DFF_529(CK,G21778,G1168);
  dff DFF_530(CK,G21779,G1169);
  dff DFF_531(CK,G21780,G1170);
  dff DFF_532(CK,G21781,G1171);
  dff DFF_533(CK,G21782,G1172);
  dff DFF_534(CK,G21783,G1173);
  dff DFF_535(CK,G21784,G1174);
  dff DFF_536(CK,G21785,G1175);
  dff DFF_537(CK,G21786,G1176);
  dff DFF_538(CK,G21787,G1177);
  dff DFF_539(CK,G21788,G1178);
  dff DFF_540(CK,G21789,G1179);
  dff DFF_541(CK,G21790,G1180);
  dff DFF_542(CK,G21791,G1181);
  dff DFF_543(CK,G21792,G1182);
  dff DFF_544(CK,G21793,G1183);
  dff DFF_545(CK,G21794,G1747);
  dff DFF_546(CK,G21795,G1184);
  dff DFF_547(CK,G21796,G1185);
  dff DFF_548(CK,G21797,G1186);
  dff DFF_549(CK,G21798,G1748);
  dff DFF_550(CK,G21799,G1187);
  dff DFF_551(CK,G21800,G1749);
  dff DFF_552(CK,G21801,G1188);
  dff DFF_553(CK,G21802,G1189);
  dff DFF_554(CK,G21803,G1750);
  dff DFF_555(CK,G21804,G1751);
  not GNAME556(G556,G1757);
  not GNAME557(G557,G1756);
  nor GNAME558(G558,G21795,G7289);
  nor GNAME559(G559,G21795,G1213);
  nand GNAME560(G560,G2010,G2011,G2012,G2013);
  nand GNAME561(G561,G2014,G2015,G2016,G2017);
  nand GNAME562(G562,G2018,G2019,G2020,G2021);
  nand GNAME563(G563,G2022,G2023,G2024,G2025);
  nand GNAME564(G564,G2026,G2027,G2028,G2029);
  nand GNAME565(G565,G2030,G2031,G2032,G2033);
  nand GNAME566(G566,G2034,G2035,G2036,G2037);
  nand GNAME567(G567,G2038,G2039,G2040,G2041);
  nand GNAME568(G568,G2042,G2043,G2044,G2045);
  nand GNAME569(G569,G2046,G2047,G2048,G2049);
  nand GNAME570(G570,G2050,G2051,G2052,G2053);
  nand GNAME571(G571,G2054,G2055,G2056,G2057);
  nand GNAME572(G572,G2058,G2059,G2060,G2061);
  nand GNAME573(G573,G2062,G2063,G2064,G2065);
  nand GNAME574(G574,G2066,G2067,G2068,G2069);
  nand GNAME575(G575,G2070,G2071,G2072,G2073);
  nand GNAME576(G576,G6736,G1272);
  nand GNAME577(G577,G6724,G6726);
  or GNAME578(G578,G2296,G577);
  nand GNAME579(G579,G6726,G1724,G6725);
  nand GNAME580(G580,G1725,G6727,G6728);
  nand GNAME581(G581,G1725,G6729,G6730);
  nand GNAME582(G582,G1725,G6731,G6732);
  nand GNAME583(G583,G1725,G6733,G6734);
  and GNAME584(G584,G5942,G2296);
  and GNAME585(G585,G5997,G2296);
  and GNAME586(G586,G6052,G2296);
  nand GNAME587(G587,G6709,G6710);
  nand GNAME588(G588,G6711,G6712);
  nand GNAME589(G589,G2295,G6713,G6714,G6715);
  nand GNAME590(G590,G7285,G7286,G1272,G6717);
  nand GNAME591(G591,G7287,G7288,G1272,G6720);
  nand GNAME592(G592,G6563,G6564,G6565,G6566);
  nand GNAME593(G593,G6570,G6571,G6569,G6567,G6568);
  nand GNAME594(G594,G6585,G6586,G6584,G6582,G6583);
  nand GNAME595(G595,G6590,G6591,G6589,G6587,G6588);
  nand GNAME596(G596,G6595,G6596,G6594,G6592,G6593);
  nand GNAME597(G597,G6600,G6601,G6599,G6597,G6598);
  nand GNAME598(G598,G6605,G6606,G6604,G6602,G6603);
  nand GNAME599(G599,G6610,G6611,G6609,G6607,G6608);
  nand GNAME600(G600,G6615,G6616,G6614,G6612,G6613);
  nand GNAME601(G601,G6620,G6621,G6619,G6617,G6618);
  nand GNAME602(G602,G6625,G6626,G6624,G6622,G6623);
  nand GNAME603(G603,G6630,G6631,G6629,G6627,G6628);
  nand GNAME604(G604,G6644,G6645,G6643,G6641,G6642);
  nand GNAME605(G605,G6649,G6650,G6648,G6646,G6647);
  nand GNAME606(G606,G6654,G6655,G6653,G6651,G6652);
  nand GNAME607(G607,G6659,G6660,G6658,G6656,G6657);
  nand GNAME608(G608,G6664,G6665,G6663,G6661,G6662);
  nand GNAME609(G609,G6669,G6670,G6668,G6666,G6667);
  nand GNAME610(G610,G6674,G6675,G6673,G6671,G6672);
  nand GNAME611(G611,G6679,G6680,G6678,G6676,G6677);
  nand GNAME612(G612,G6684,G6685,G6683,G6681,G6682);
  nand GNAME613(G613,G6689,G6690,G6688,G6686,G6687);
  nand GNAME614(G614,G6536,G6537,G6535,G6533,G6534);
  nand GNAME615(G615,G6541,G6542,G6540,G6538,G6539);
  nand GNAME616(G616,G6546,G6547,G6545,G6543,G6544);
  nand GNAME617(G617,G6551,G6552,G6550,G6548,G6549);
  nand GNAME618(G618,G6556,G6557,G6555,G6553,G6554);
  nand GNAME619(G619,G6561,G6562,G6560,G6558,G6559);
  nand GNAME620(G620,G2244,G6578,G6579,G6580,G6581);
  nand GNAME621(G621,G2245,G6637,G6638,G6639,G6640);
  nand GNAME622(G622,G2246,G6691,G6693,G6698,G6699);
  nand GNAME623(G623,G2247,G6700,G6702,G6707,G6708);
  and GNAME624(G624,G568,G1571);
  and GNAME625(G625,G569,G1571);
  and GNAME626(G626,G570,G1571);
  and GNAME627(G627,G571,G1571);
  and GNAME628(G628,G572,G1571);
  and GNAME629(G629,G573,G1571);
  and GNAME630(G630,G574,G1571);
  and GNAME631(G631,G575,G1571);
  nand GNAME632(G632,G1558,G1715,G2301,G2298,G1713);
  nand GNAME633(G633,G1713,G2317,G6530,G1722);
  nand GNAME634(G634,G6405,G6406,G6407,G6408);
  nand GNAME635(G635,G6412,G6413,G6411,G6409,G6410);
  nand GNAME636(G636,G6427,G6428,G6426,G6424,G6425);
  nand GNAME637(G637,G6432,G6433,G6431,G6429,G6430);
  nand GNAME638(G638,G6437,G6438,G6436,G6434,G6435);
  nand GNAME639(G639,G6442,G6443,G6441,G6439,G6440);
  nand GNAME640(G640,G6447,G6448,G6446,G6444,G6445);
  nand GNAME641(G641,G6452,G6453,G6451,G6449,G6450);
  nand GNAME642(G642,G6457,G6458,G6456,G6454,G6455);
  nand GNAME643(G643,G6459,G6460,G6461,G6462);
  nand GNAME644(G644,G6463,G6464,G6465,G6466);
  nand GNAME645(G645,G6467,G6468,G6469,G6470);
  nand GNAME646(G646,G6476,G6477,G6478,G6479);
  nand GNAME647(G647,G6480,G6481,G6482,G6483);
  nand GNAME648(G648,G6484,G6485,G6486,G6487);
  nand GNAME649(G649,G6488,G6489,G6490,G6491);
  nand GNAME650(G650,G6492,G6493,G6494,G6495);
  nand GNAME651(G651,G6496,G6497,G6498,G6499);
  nand GNAME652(G652,G6500,G6501,G6502,G6503);
  nand GNAME653(G653,G6504,G6505,G6506,G6507);
  nand GNAME654(G654,G6508,G6509,G6510,G6511);
  nand GNAME655(G655,G6512,G6513,G6514,G6515);
  nand GNAME656(G656,G6379,G6380,G6381,G6382);
  nand GNAME657(G657,G6383,G6384,G6385,G6386);
  nand GNAME658(G658,G6387,G6388,G6389,G6390);
  nand GNAME659(G659,G6391,G6392,G6393,G6394);
  nand GNAME660(G660,G6395,G6396,G6397,G6398);
  nand GNAME661(G661,G6403,G6404,G6402,G6400,G6401);
  nand GNAME662(G662,G6422,G6423,G6421,G6419,G6420);
  nand GNAME663(G663,G6474,G6475,G6473,G6471,G6472);
  nand GNAME664(G664,G6519,G6520,G6518,G6516,G6517);
  nand GNAME665(G665,G6524,G6525,G6523,G6521,G6522);
  and GNAME666(G666,G5959,G2300);
  and GNAME667(G667,G6014,G2300);
  and GNAME668(G668,G6069,G2300);
  and GNAME669(G669,G6124,G2300);
  and GNAME670(G670,G6180,G2300);
  and GNAME671(G671,G6236,G2300);
  and GNAME672(G672,G6292,G2300);
  and GNAME673(G673,G6348,G2300);
  and GNAME674(G674,G21549,G1571);
  and GNAME675(G675,G21550,G1571);
  and GNAME676(G676,G21551,G1571);
  and GNAME677(G677,G21552,G1571);
  and GNAME678(G678,G21553,G1571);
  nand GNAME679(G679,G6354,G2305,G2307);
  nand GNAME680(G680,G1715,G2238,G2306,G1551,G2304);
  nand GNAME681(G681,G2305,G2317,G6363,G6364);
  and GNAME682(G682,G1242,G2545);
  and GNAME683(G683,G1238,G2477);
  or GNAME684(G684,G21567,G7296);
  nand GNAME685(G685,G5960,G5961,G5962,G5963);
  nand GNAME686(G686,G6015,G6016,G6017,G6018);
  nand GNAME687(G687,G6070,G6071,G6072,G6073);
  nand GNAME688(G688,G6128,G6129,G6127,G6125,G6126);
  nand GNAME689(G689,G6184,G6185,G6183,G6181,G6182);
  nand GNAME690(G690,G2211,G6238,G6239,G6240);
  nand GNAME691(G691,G2224,G6294,G6295,G6296);
  nand GNAME692(G692,G2237,G6350,G6351,G6352);
  nand GNAME693(G693,G5780,G5781,G5782,G5783);
  nand GNAME694(G694,G5787,G5788,G5786,G5784,G5785);
  nand GNAME695(G695,G5797,G5798,G5796,G5794,G5795);
  nand GNAME696(G696,G5802,G5803,G5801,G5799,G5800);
  nand GNAME697(G697,G5807,G5808,G5806,G5804,G5805);
  nand GNAME698(G698,G5812,G5813,G5811,G5809,G5810);
  nand GNAME699(G699,G5817,G5818,G5816,G5814,G5815);
  nand GNAME700(G700,G5822,G5823,G5821,G5819,G5820);
  nand GNAME701(G701,G5827,G5828,G5826,G5824,G5825);
  nand GNAME702(G702,G5832,G5833,G5831,G5829,G5830);
  nand GNAME703(G703,G5837,G5838,G5836,G5834,G5835);
  nand GNAME704(G704,G5842,G5843,G5841,G5839,G5840);
  nand GNAME705(G705,G5852,G5853,G5851,G5849,G5850);
  nand GNAME706(G706,G5857,G5858,G5856,G5854,G5855);
  nand GNAME707(G707,G5862,G5863,G5861,G5859,G5860);
  nand GNAME708(G708,G5867,G5868,G5866,G5864,G5865);
  nand GNAME709(G709,G5872,G5873,G5871,G5869,G5870);
  nand GNAME710(G710,G5877,G5878,G5876,G5874,G5875);
  nand GNAME711(G711,G5882,G5883,G5881,G5879,G5880);
  nand GNAME712(G712,G5887,G5888,G5886,G5884,G5885);
  nand GNAME713(G713,G5892,G5893,G5891,G5889,G5890);
  nand GNAME714(G714,G5897,G5898,G5896,G5894,G5895);
  nand GNAME715(G715,G5753,G5754,G5752,G5750,G5751);
  nand GNAME716(G716,G5758,G5759,G5757,G5755,G5756);
  nand GNAME717(G717,G5763,G5764,G5762,G5760,G5761);
  nand GNAME718(G718,G5768,G5769,G5767,G5765,G5766);
  nand GNAME719(G719,G5773,G5774,G5772,G5770,G5771);
  nand GNAME720(G720,G5778,G5779,G5777,G5775,G5776);
  nand GNAME721(G721,G5792,G5793,G5791,G5789,G5790);
  nand GNAME722(G722,G5847,G5848,G5846,G5844,G5845);
  nand GNAME723(G723,G5902,G5903,G5901,G5899,G5900);
  nand GNAME724(G724,G2138,G5906,G5904,G5905);
  and GNAME725(G725,G2511,G21598);
  and GNAME726(G726,G2511,G21589);
  and GNAME727(G727,G2511,G21588);
  and GNAME728(G728,G2511,G21587);
  and GNAME729(G729,G2511,G21586);
  and GNAME730(G730,G2511,G21585);
  and GNAME731(G731,G2511,G21584);
  and GNAME732(G732,G2511,G21583);
  and GNAME733(G733,G2511,G21582);
  and GNAME734(G734,G2511,G21581);
  and GNAME735(G735,G2511,G21580);
  and GNAME736(G736,G2511,G21579);
  and GNAME737(G737,G2511,G21578);
  and GNAME738(G738,G2511,G21577);
  and GNAME739(G739,G2511,G21576);
  and GNAME740(G740,G2511,G21575);
  and GNAME741(G741,G2511,G21574);
  and GNAME742(G742,G2511,G21573);
  and GNAME743(G743,G2511,G21572);
  and GNAME744(G744,G2511,G21571);
  and GNAME745(G745,G2511,G21570);
  and GNAME746(G746,G2511,G21569);
  and GNAME747(G747,G2511,G21568);
  and GNAME748(G748,G2511,G21567);
  and GNAME749(G749,G1248,G5492);
  and GNAME750(G750,G1248,G5509);
  and GNAME751(G751,G1248,G5526);
  and GNAME752(G752,G1248,G5543);
  and GNAME753(G753,G1248,G5560);
  and GNAME754(G754,G1248,G5577);
  and GNAME755(G755,G1248,G5594);
  and GNAME756(G756,G1248,G5611);
  nand GNAME757(G757,G2353,G2351,G2352);
  nand GNAME758(G758,G2356,G2354,G2355);
  nand GNAME759(G759,G2359,G2357,G2358);
  nand GNAME760(G760,G2362,G2360,G2361);
  nand GNAME761(G761,G2365,G2363,G2364);
  nand GNAME762(G762,G2368,G2366,G2367);
  nand GNAME763(G763,G2371,G2369,G2370);
  nand GNAME764(G764,G2374,G2372,G2373);
  nand GNAME765(G765,G2377,G2375,G2376);
  nand GNAME766(G766,G2380,G2378,G2379);
  nand GNAME767(G767,G2383,G2381,G2382);
  nand GNAME768(G768,G2386,G2384,G2385);
  nand GNAME769(G769,G2389,G2387,G2388);
  nand GNAME770(G770,G2392,G2390,G2391);
  nand GNAME771(G771,G2395,G2393,G2394);
  nand GNAME772(G772,G2398,G2396,G2397);
  nand GNAME773(G773,G2401,G2399,G2400);
  nand GNAME774(G774,G2404,G2402,G2403);
  nand GNAME775(G775,G2407,G2405,G2406);
  nand GNAME776(G776,G2410,G2408,G2409);
  nand GNAME777(G777,G2413,G2411,G2412);
  nand GNAME778(G778,G2416,G2414,G2415);
  nand GNAME779(G779,G2419,G2417,G2418);
  nand GNAME780(G780,G2422,G2420,G2421);
  nand GNAME781(G781,G2425,G2423,G2424);
  nand GNAME782(G782,G2428,G2426,G2427);
  nand GNAME783(G783,G2431,G2429,G2430);
  nand GNAME784(G784,G2434,G2432,G2433);
  nand GNAME785(G785,G2437,G2435,G2436);
  nand GNAME786(G786,G2440,G2438,G2439);
  nand GNAME787(G787,G2449,G2335,G2448);
  or GNAME788(G788,G36,G7292);
  nand GNAME789(G789,G6766,G6767,G2336,G2452);
  or GNAME790(G790,G6768,G6769,G1203,G1200);
  and GNAME791(G791,G6772,G21395);
  and GNAME792(G792,G6772,G21396);
  and GNAME793(G793,G6772,G21397);
  and GNAME794(G794,G6772,G21398);
  and GNAME795(G795,G6772,G21399);
  and GNAME796(G796,G6772,G21400);
  and GNAME797(G797,G6772,G21401);
  and GNAME798(G798,G6772,G21402);
  and GNAME799(G799,G6772,G21403);
  and GNAME800(G800,G6772,G21404);
  and GNAME801(G801,G6772,G21405);
  and GNAME802(G802,G6772,G21406);
  and GNAME803(G803,G6772,G21407);
  and GNAME804(G804,G6772,G21408);
  and GNAME805(G805,G6772,G21409);
  and GNAME806(G806,G6772,G21410);
  and GNAME807(G807,G6772,G21411);
  and GNAME808(G808,G6772,G21412);
  and GNAME809(G809,G6772,G21413);
  and GNAME810(G810,G6772,G21414);
  and GNAME811(G811,G6772,G21415);
  and GNAME812(G812,G6772,G21416);
  and GNAME813(G813,G6772,G21417);
  and GNAME814(G814,G6772,G21418);
  and GNAME815(G815,G6772,G21419);
  and GNAME816(G816,G6772,G21420);
  and GNAME817(G817,G6772,G21421);
  and GNAME818(G818,G6772,G21422);
  and GNAME819(G819,G6772,G21423);
  and GNAME820(G820,G6772,G21424);
  or GNAME821(G821,G1274,G1291,G6749);
  nand GNAME822(G822,G2306,G2332,G2616,G2617);
  nand GNAME823(G823,G2622,G2342,G2621);
  nand GNAME824(G824,G6779,G6780,G2341,G2343);
  nand GNAME825(G825,G1804,G2703,G2701,G2702);
  nand GNAME826(G826,G1805,G2716,G2714,G2715);
  nand GNAME827(G827,G1806,G2729,G2727,G2728);
  nand GNAME828(G828,G1807,G2742,G2740,G2741);
  nand GNAME829(G829,G1808,G2755,G2753,G2754);
  nand GNAME830(G830,G1809,G2768,G2766,G2767);
  nand GNAME831(G831,G1810,G2781,G2779,G2780);
  nand GNAME832(G832,G1811,G2794,G2792,G2793);
  nand GNAME833(G833,G1812,G2811,G2809,G2810);
  nand GNAME834(G834,G1813,G2821,G2819,G2820);
  nand GNAME835(G835,G1814,G2831,G2829,G2830);
  nand GNAME836(G836,G1815,G2841,G2839,G2840);
  nand GNAME837(G837,G1816,G2851,G2849,G2850);
  nand GNAME838(G838,G1817,G2861,G2859,G2860);
  nand GNAME839(G839,G1818,G2871,G2869,G2870);
  nand GNAME840(G840,G1819,G2881,G2879,G2880);
  nand GNAME841(G841,G1820,G2898,G2896,G2897);
  nand GNAME842(G842,G1821,G2908,G2906,G2907);
  nand GNAME843(G843,G1822,G2918,G2916,G2917);
  nand GNAME844(G844,G1823,G2928,G2926,G2927);
  nand GNAME845(G845,G1824,G2938,G2936,G2937);
  nand GNAME846(G846,G1825,G2948,G2946,G2947);
  nand GNAME847(G847,G1826,G2958,G2956,G2957);
  nand GNAME848(G848,G1827,G2968,G2966,G2967);
  nand GNAME849(G849,G1828,G2985,G2983,G2984);
  nand GNAME850(G850,G1829,G2995,G2993,G2994);
  nand GNAME851(G851,G1830,G3005,G3003,G3004);
  nand GNAME852(G852,G1831,G3015,G3013,G3014);
  nand GNAME853(G853,G1832,G3025,G3023,G3024);
  nand GNAME854(G854,G1833,G3035,G3033,G3034);
  nand GNAME855(G855,G1834,G3045,G3043,G3044);
  nand GNAME856(G856,G1835,G3055,G3053,G3054);
  nand GNAME857(G857,G1836,G3072,G3070,G3071);
  nand GNAME858(G858,G1837,G3082,G3080,G3081);
  nand GNAME859(G859,G1838,G3092,G3090,G3091);
  nand GNAME860(G860,G1839,G3102,G3100,G3101);
  nand GNAME861(G861,G1840,G3112,G3110,G3111);
  nand GNAME862(G862,G1841,G3122,G3120,G3121);
  nand GNAME863(G863,G1842,G3132,G3130,G3131);
  nand GNAME864(G864,G1843,G3142,G3140,G3141);
  nand GNAME865(G865,G1844,G3159,G3157,G3158);
  nand GNAME866(G866,G1845,G3169,G3167,G3168);
  nand GNAME867(G867,G1846,G3179,G3177,G3178);
  nand GNAME868(G868,G1847,G3189,G3187,G3188);
  nand GNAME869(G869,G1848,G3199,G3197,G3198);
  nand GNAME870(G870,G1849,G3209,G3207,G3208);
  nand GNAME871(G871,G1850,G3219,G3217,G3218);
  nand GNAME872(G872,G1851,G3229,G3227,G3228);
  nand GNAME873(G873,G1852,G3246,G3244,G3245);
  nand GNAME874(G874,G1853,G3256,G3254,G3255);
  nand GNAME875(G875,G1854,G3266,G3264,G3265);
  nand GNAME876(G876,G1855,G3276,G3274,G3275);
  nand GNAME877(G877,G1856,G3286,G3284,G3285);
  nand GNAME878(G878,G1857,G3296,G3294,G3295);
  nand GNAME879(G879,G1858,G3306,G3304,G3305);
  nand GNAME880(G880,G1859,G3316,G3314,G3315);
  nand GNAME881(G881,G1860,G3333,G3331,G3332);
  nand GNAME882(G882,G1861,G3343,G3341,G3342);
  nand GNAME883(G883,G1862,G3353,G3351,G3352);
  nand GNAME884(G884,G1863,G3363,G3361,G3362);
  nand GNAME885(G885,G1864,G3373,G3371,G3372);
  nand GNAME886(G886,G1865,G3383,G3381,G3382);
  nand GNAME887(G887,G1866,G3393,G3391,G3392);
  nand GNAME888(G888,G1867,G3403,G3401,G3402);
  nand GNAME889(G889,G1868,G3420,G3418,G3419);
  nand GNAME890(G890,G1869,G3430,G3428,G3429);
  nand GNAME891(G891,G1870,G3440,G3438,G3439);
  nand GNAME892(G892,G1871,G3450,G3448,G3449);
  nand GNAME893(G893,G1872,G3460,G3458,G3459);
  nand GNAME894(G894,G1873,G3470,G3468,G3469);
  nand GNAME895(G895,G1874,G3480,G3478,G3479);
  nand GNAME896(G896,G1875,G3490,G3488,G3489);
  nand GNAME897(G897,G1876,G3507,G3505,G3506);
  nand GNAME898(G898,G1877,G3517,G3515,G3516);
  nand GNAME899(G899,G1878,G3527,G3525,G3526);
  nand GNAME900(G900,G1879,G3537,G3535,G3536);
  nand GNAME901(G901,G1880,G3547,G3545,G3546);
  nand GNAME902(G902,G1881,G3557,G3555,G3556);
  nand GNAME903(G903,G1882,G3567,G3565,G3566);
  nand GNAME904(G904,G1883,G3577,G3575,G3576);
  nand GNAME905(G905,G1884,G3594,G3592,G3593);
  nand GNAME906(G906,G1885,G3604,G3602,G3603);
  nand GNAME907(G907,G1886,G3614,G3612,G3613);
  nand GNAME908(G908,G1887,G3624,G3622,G3623);
  nand GNAME909(G909,G1888,G3634,G3632,G3633);
  nand GNAME910(G910,G1889,G3644,G3642,G3643);
  nand GNAME911(G911,G1890,G3654,G3652,G3653);
  nand GNAME912(G912,G1891,G3664,G3662,G3663);
  nand GNAME913(G913,G1892,G3681,G3679,G3680);
  nand GNAME914(G914,G1893,G3691,G3689,G3690);
  nand GNAME915(G915,G1894,G3701,G3699,G3700);
  nand GNAME916(G916,G1895,G3711,G3709,G3710);
  nand GNAME917(G917,G1896,G3721,G3719,G3720);
  nand GNAME918(G918,G1897,G3731,G3729,G3730);
  nand GNAME919(G919,G1898,G3741,G3739,G3740);
  nand GNAME920(G920,G1899,G3751,G3749,G3750);
  nand GNAME921(G921,G1900,G3768,G3766,G3767);
  nand GNAME922(G922,G1901,G3778,G3776,G3777);
  nand GNAME923(G923,G1902,G3788,G3786,G3787);
  nand GNAME924(G924,G1903,G3798,G3796,G3797);
  nand GNAME925(G925,G1904,G3808,G3806,G3807);
  nand GNAME926(G926,G1905,G3818,G3816,G3817);
  nand GNAME927(G927,G1906,G3828,G3826,G3827);
  nand GNAME928(G928,G1907,G3838,G3836,G3837);
  nand GNAME929(G929,G1908,G3855,G3853,G3854);
  nand GNAME930(G930,G1909,G3865,G3863,G3864);
  nand GNAME931(G931,G1910,G3875,G3873,G3874);
  nand GNAME932(G932,G1911,G3885,G3883,G3884);
  nand GNAME933(G933,G1912,G3895,G3893,G3894);
  nand GNAME934(G934,G1913,G3905,G3903,G3904);
  nand GNAME935(G935,G1914,G3915,G3913,G3914);
  nand GNAME936(G936,G1915,G3925,G3923,G3924);
  nand GNAME937(G937,G1916,G3942,G3940,G3941);
  nand GNAME938(G938,G1917,G3952,G3950,G3951);
  nand GNAME939(G939,G1918,G3962,G3960,G3961);
  nand GNAME940(G940,G1919,G3972,G3970,G3971);
  nand GNAME941(G941,G1920,G3982,G3980,G3981);
  nand GNAME942(G942,G1921,G3992,G3990,G3991);
  nand GNAME943(G943,G1922,G4002,G4000,G4001);
  nand GNAME944(G944,G1923,G4012,G4010,G4011);
  nand GNAME945(G945,G1924,G4029,G4027,G4028);
  nand GNAME946(G946,G1925,G4039,G4037,G4038);
  nand GNAME947(G947,G1926,G4049,G4047,G4048);
  nand GNAME948(G948,G1927,G4059,G4057,G4058);
  nand GNAME949(G949,G1928,G4069,G4067,G4068);
  nand GNAME950(G950,G1929,G4079,G4077,G4078);
  nand GNAME951(G951,G1930,G4089,G4087,G4088);
  nand GNAME952(G952,G1931,G4099,G4097,G4098);
  nor GNAME953(G953,G1532,G7293);
  nand GNAME954(G954,G4189,G4187,G4188);
  nand GNAME955(G955,G4192,G4190,G4191);
  nand GNAME956(G956,G4195,G4193,G4194);
  nand GNAME957(G957,G1938,G4213,G4216,G4217);
  nand GNAME958(G958,G1939,G4219,G4222,G4223);
  nand GNAME959(G959,G1940,G4225,G4228,G4229);
  nand GNAME960(G960,G1941,G4231,G4234,G4235);
  nand GNAME961(G961,G1942,G4237,G4240,G4241);
  nand GNAME962(G962,G1943,G4243,G4246,G4247);
  nand GNAME963(G963,G1944,G4249,G4252,G4253);
  nand GNAME964(G964,G1945,G4255,G4258,G4259);
  nand GNAME965(G965,G1946,G4261,G4264,G4265);
  nand GNAME966(G966,G1947,G4267,G4270,G4271);
  nand GNAME967(G967,G1948,G4273,G4276,G4277);
  nand GNAME968(G968,G1949,G4279,G4282,G4283);
  nand GNAME969(G969,G1950,G4285,G4288,G4289);
  nand GNAME970(G970,G1951,G4291,G4294,G4295);
  nand GNAME971(G971,G1952,G4297,G4300,G4301);
  nand GNAME972(G972,G1953,G4303,G4306,G4307);
  nand GNAME973(G973,G1954,G4309,G4312,G4313);
  nand GNAME974(G974,G1955,G4315,G4318,G4319);
  nand GNAME975(G975,G1956,G4321,G4324,G4325);
  nand GNAME976(G976,G1957,G4327,G4330,G4331);
  nand GNAME977(G977,G1958,G4333,G4336,G4337);
  nand GNAME978(G978,G1959,G4339,G4342,G4343);
  nand GNAME979(G979,G1960,G4345,G4348,G4349);
  nand GNAME980(G980,G1961,G4351,G4354,G4355);
  nand GNAME981(G981,G1962,G4357,G4360,G4361);
  nand GNAME982(G982,G1963,G4363,G4366,G4367);
  nand GNAME983(G983,G1964,G4369,G4372,G4373);
  nand GNAME984(G984,G1965,G4375,G4378,G4379);
  nand GNAME985(G985,G1966,G4381,G4384,G4385);
  nand GNAME986(G986,G1967,G4387,G4390,G4391);
  nand GNAME987(G987,G1968,G4393,G4396,G4397);
  nand GNAME988(G988,G1969,G4399,G4402,G4403);
  nand GNAME989(G989,G4410,G4411,G4409,G4407,G4408);
  nand GNAME990(G990,G4415,G4416,G4414,G4412,G4413);
  nand GNAME991(G991,G4420,G4421,G4419,G4417,G4418);
  nand GNAME992(G992,G4425,G4426,G4424,G4422,G4423);
  nand GNAME993(G993,G4430,G4431,G4429,G4427,G4428);
  nand GNAME994(G994,G4435,G4436,G4434,G4432,G4433);
  nand GNAME995(G995,G4440,G4441,G4439,G4437,G4438);
  nand GNAME996(G996,G4445,G4446,G4444,G4442,G4443);
  nand GNAME997(G997,G4450,G4451,G4449,G4447,G4448);
  nand GNAME998(G998,G4455,G4456,G4454,G4452,G4453);
  nand GNAME999(G999,G4460,G4461,G4459,G4457,G4458);
  nand GNAME1000(G1000,G4465,G4466,G4464,G4462,G4463);
  nand GNAME1001(G1001,G4470,G4471,G4469,G4467,G4468);
  nand GNAME1002(G1002,G4475,G4476,G4474,G4472,G4473);
  nand GNAME1003(G1003,G4480,G4481,G4479,G4477,G4478);
  nand GNAME1004(G1004,G4485,G4486,G4484,G4482,G4483);
  nand GNAME1005(G1005,G4490,G4491,G4489,G4487,G4488);
  nand GNAME1006(G1006,G4495,G4496,G4494,G4492,G4493);
  nand GNAME1007(G1007,G4500,G4501,G4499,G4497,G4498);
  nand GNAME1008(G1008,G4505,G4506,G4504,G4502,G4503);
  nand GNAME1009(G1009,G4510,G4511,G4509,G4507,G4508);
  nand GNAME1010(G1010,G4515,G4516,G4514,G4512,G4513);
  nand GNAME1011(G1011,G4520,G4521,G4519,G4517,G4518);
  nand GNAME1012(G1012,G4525,G4526,G4524,G4522,G4523);
  nand GNAME1013(G1013,G4530,G4531,G4529,G4527,G4528);
  nand GNAME1014(G1014,G4535,G4536,G4534,G4532,G4533);
  nand GNAME1015(G1015,G4540,G4541,G4539,G4537,G4538);
  nand GNAME1016(G1016,G4545,G4546,G4544,G4542,G4543);
  nand GNAME1017(G1017,G4550,G4551,G4549,G4547,G4548);
  nand GNAME1018(G1018,G4555,G4556,G4554,G4552,G4553);
  nand GNAME1019(G1019,G4560,G4561,G4559,G4557,G4558);
  nand GNAME1020(G1020,G4565,G4566,G4564,G4562,G4563);
  nand GNAME1021(G1021,G4571,G4569,G4570);
  nand GNAME1022(G1022,G4573,G4572,G4603);
  nand GNAME1023(G1023,G4575,G4574,G4606);
  nand GNAME1024(G1024,G4577,G4576,G4609);
  nand GNAME1025(G1025,G4579,G4578,G4612);
  nand GNAME1026(G1026,G4581,G4580,G4615);
  nand GNAME1027(G1027,G4583,G4582,G4618);
  nand GNAME1028(G1028,G4585,G4584,G4621);
  nand GNAME1029(G1029,G4587,G4586,G4624);
  nand GNAME1030(G1030,G4589,G4588,G4627);
  nand GNAME1031(G1031,G4591,G4590,G4630);
  nand GNAME1032(G1032,G4593,G4592,G4633);
  nand GNAME1033(G1033,G4595,G4594,G4636);
  nand GNAME1034(G1034,G4597,G4596,G4639);
  nand GNAME1035(G1035,G4599,G4598,G4642);
  nand GNAME1036(G1036,G4601,G4600,G4645);
  nand GNAME1037(G1037,G4604,G4602,G4603);
  nand GNAME1038(G1038,G4607,G4605,G4606);
  nand GNAME1039(G1039,G4610,G4608,G4609);
  nand GNAME1040(G1040,G4613,G4611,G4612);
  nand GNAME1041(G1041,G4616,G4614,G4615);
  nand GNAME1042(G1042,G4619,G4617,G4618);
  nand GNAME1043(G1043,G4622,G4620,G4621);
  nand GNAME1044(G1044,G4625,G4623,G4624);
  nand GNAME1045(G1045,G4628,G4626,G4627);
  nand GNAME1046(G1046,G4631,G4629,G4630);
  nand GNAME1047(G1047,G4634,G4632,G4633);
  nand GNAME1048(G1048,G4637,G4635,G4636);
  nand GNAME1049(G1049,G4640,G4638,G4639);
  nand GNAME1050(G1050,G4643,G4641,G4642);
  nand GNAME1051(G1051,G4646,G4644,G4645);
  nand GNAME1052(G1052,G4654,G4652,G4653);
  nand GNAME1053(G1053,G4657,G4655,G4656);
  nand GNAME1054(G1054,G4660,G4658,G4659);
  nand GNAME1055(G1055,G4663,G4661,G4662);
  nand GNAME1056(G1056,G4666,G4664,G4665);
  nand GNAME1057(G1057,G4669,G4667,G4668);
  nand GNAME1058(G1058,G4672,G4670,G4671);
  nand GNAME1059(G1059,G4675,G4673,G4674);
  nand GNAME1060(G1060,G4678,G4676,G4677);
  nand GNAME1061(G1061,G4681,G4679,G4680);
  nand GNAME1062(G1062,G4684,G4682,G4683);
  nand GNAME1063(G1063,G4687,G4685,G4686);
  nand GNAME1064(G1064,G4690,G4688,G4689);
  nand GNAME1065(G1065,G4693,G4691,G4692);
  nand GNAME1066(G1066,G4696,G4694,G4695);
  nand GNAME1067(G1067,G4699,G4697,G4698);
  nand GNAME1068(G1068,G4702,G4700,G4701);
  nand GNAME1069(G1069,G4705,G4703,G4704);
  nand GNAME1070(G1070,G4708,G4706,G4707);
  nand GNAME1071(G1071,G4711,G4709,G4710);
  nand GNAME1072(G1072,G4714,G4712,G4713);
  nand GNAME1073(G1073,G4717,G4715,G4716);
  nand GNAME1074(G1074,G4720,G4718,G4719);
  nand GNAME1075(G1075,G4723,G4721,G4722);
  nand GNAME1076(G1076,G4726,G4724,G4725);
  nand GNAME1077(G1077,G4729,G4727,G4728);
  nand GNAME1078(G1078,G4732,G4730,G4731);
  nand GNAME1079(G1079,G4735,G4733,G4734);
  nand GNAME1080(G1080,G4738,G4736,G4737);
  nand GNAME1081(G1081,G4741,G4739,G4740);
  nand GNAME1082(G1082,G4744,G4742,G4743);
  and GNAME1083(G1083,G1561,G21693);
  nand GNAME1084(G1084,G4749,G4750,G4751,G4752);
  nand GNAME1085(G1085,G4753,G4754,G4755,G4756);
  nand GNAME1086(G1086,G4757,G4758,G4759,G4760);
  nand GNAME1087(G1087,G4761,G4762,G4763,G4764);
  nand GNAME1088(G1088,G4765,G4766,G4767,G4768);
  nand GNAME1089(G1089,G4769,G4770,G4771,G4772);
  nand GNAME1090(G1090,G4773,G4774,G4775,G4776);
  nand GNAME1091(G1091,G4777,G4778,G4779,G4780);
  nand GNAME1092(G1092,G4781,G4782,G4783,G4784);
  nand GNAME1093(G1093,G4785,G4786,G4787,G4788);
  nand GNAME1094(G1094,G4789,G4790,G4791,G4792);
  nand GNAME1095(G1095,G4793,G4794,G4795,G4796);
  nand GNAME1096(G1096,G4797,G4798,G4799,G4800);
  nand GNAME1097(G1097,G4801,G4802,G4803,G4804);
  nand GNAME1098(G1098,G4805,G4806,G4807,G4808);
  nand GNAME1099(G1099,G4809,G4810,G4811,G4812);
  nand GNAME1100(G1100,G4816,G4817,G4815,G4813,G4814);
  nand GNAME1101(G1101,G4821,G4822,G4820,G4818,G4819);
  nand GNAME1102(G1102,G4826,G4827,G4825,G4823,G4824);
  nand GNAME1103(G1103,G4831,G4832,G4830,G4828,G4829);
  nand GNAME1104(G1104,G4836,G4837,G4835,G4833,G4834);
  nand GNAME1105(G1105,G4841,G4842,G4840,G4838,G4839);
  nand GNAME1106(G1106,G4846,G4847,G4845,G4843,G4844);
  nand GNAME1107(G1107,G4851,G4852,G4850,G4848,G4849);
  nand GNAME1108(G1108,G4856,G4857,G4855,G4853,G4854);
  nand GNAME1109(G1109,G4861,G4862,G4860,G4858,G4859);
  nand GNAME1110(G1110,G4866,G4867,G4865,G4863,G4864);
  nand GNAME1111(G1111,G4871,G4872,G4870,G4868,G4869);
  nand GNAME1112(G1112,G4876,G4877,G4875,G4873,G4874);
  nand GNAME1113(G1113,G4881,G4882,G4880,G4878,G4879);
  nand GNAME1114(G1114,G4886,G4887,G4885,G4883,G4884);
  nand GNAME1115(G1115,G4890,G4888,G4889);
  nand GNAME1116(G1116,G4895,G4893,G4894);
  nand GNAME1117(G1117,G4898,G4896,G4897);
  nand GNAME1118(G1118,G4901,G4899,G4900);
  nand GNAME1119(G1119,G4904,G4902,G4903);
  nand GNAME1120(G1120,G4907,G4905,G4906);
  nand GNAME1121(G1121,G4910,G4908,G4909);
  nand GNAME1122(G1122,G4913,G4911,G4912);
  nand GNAME1123(G1123,G4916,G4914,G4915);
  nand GNAME1124(G1124,G4919,G4917,G4918);
  nand GNAME1125(G1125,G4922,G4920,G4921);
  nand GNAME1126(G1126,G4925,G4923,G4924);
  nand GNAME1127(G1127,G4928,G4926,G4927);
  nand GNAME1128(G1128,G4931,G4929,G4930);
  nand GNAME1129(G1129,G4934,G4932,G4933);
  nand GNAME1130(G1130,G4937,G4935,G4936);
  nand GNAME1131(G1131,G4940,G4938,G4939);
  nand GNAME1132(G1132,G4943,G4941,G4942);
  nand GNAME1133(G1133,G4946,G4944,G4945);
  nand GNAME1134(G1134,G4949,G4947,G4948);
  nand GNAME1135(G1135,G4952,G4950,G4951);
  nand GNAME1136(G1136,G4955,G4953,G4954);
  nand GNAME1137(G1137,G4958,G4956,G4957);
  nand GNAME1138(G1138,G4961,G4959,G4960);
  nand GNAME1139(G1139,G4964,G4962,G4963);
  nand GNAME1140(G1140,G4967,G4965,G4966);
  nand GNAME1141(G1141,G4970,G4968,G4969);
  nand GNAME1142(G1142,G4973,G4971,G4972);
  nand GNAME1143(G1143,G4976,G4974,G4975);
  nand GNAME1144(G1144,G4979,G4977,G4978);
  nand GNAME1145(G1145,G4982,G4980,G4981);
  nand GNAME1146(G1146,G4985,G4983,G4984);
  nand GNAME1147(G1147,G4986,G4987);
  nand GNAME1148(G1148,G1970,G5001,G4998,G4999);
  nand GNAME1149(G1149,G1971,G5007,G5004,G5005);
  nand GNAME1150(G1150,G1972,G5013,G5010,G5011);
  nand GNAME1151(G1151,G1973,G5019,G5016,G5017);
  nand GNAME1152(G1152,G1974,G5025,G5022,G5023,G5024);
  nand GNAME1153(G1153,G1975,G5031,G5028,G5029,G5030);
  nand GNAME1154(G1154,G1976,G5037,G5034,G5035,G5036);
  nand GNAME1155(G1155,G1977,G5043,G5040,G5041,G5042);
  nand GNAME1156(G1156,G1978,G5049,G5046,G5047,G5048);
  nand GNAME1157(G1157,G1979,G5055,G5052,G5053,G5054);
  nand GNAME1158(G1158,G1980,G5061,G5058,G5059,G5060);
  nand GNAME1159(G1159,G1981,G5067,G5064,G5065,G5066);
  nand GNAME1160(G1160,G1982,G5073,G5070,G5071,G5072);
  nand GNAME1161(G1161,G1983,G5079,G5076,G5077,G5078);
  nand GNAME1162(G1162,G1984,G5085,G5082,G5083,G5084);
  nand GNAME1163(G1163,G1985,G5091,G5088,G5089,G5090);
  nand GNAME1164(G1164,G1986,G5097,G5094,G5095,G5096);
  nand GNAME1165(G1165,G1987,G5103,G5100,G5101,G5102);
  nand GNAME1166(G1166,G1988,G5109,G5106,G5107,G5108);
  nand GNAME1167(G1167,G1989,G5115,G5112,G5113,G5114);
  nand GNAME1168(G1168,G1990,G5121,G5118,G5119);
  nand GNAME1169(G1169,G1991,G5127,G5124,G5125);
  nand GNAME1170(G1170,G1992,G5133,G5130,G5131);
  nand GNAME1171(G1171,G1993,G5139,G5136,G5137);
  nand GNAME1172(G1172,G1994,G5145,G5142,G5143);
  nand GNAME1173(G1173,G1995,G5150,G5148,G5149);
  nand GNAME1174(G1174,G1996,G5156,G5154,G5155);
  nand GNAME1175(G1175,G1997,G5162,G5160,G5161);
  nand GNAME1176(G1176,G1998,G5168,G5166,G5167);
  nand GNAME1177(G1177,G1999,G5174,G5172,G5173);
  nand GNAME1178(G1178,G2000,G5180,G5178,G5179);
  nand GNAME1179(G1179,G2001,G5186,G5184,G5185);
  nand GNAME1180(G1180,G2339,G7220,G7221);
  nand GNAME1181(G1181,G5191,G7222,G7223);
  nand GNAME1182(G1182,G5192,G2339,G1587);
  nand GNAME1183(G1183,G1587,G7224,G7225);
  nand GNAME1184(G1184,G5194,G5195);
  nand GNAME1185(G1185,G5204,G5205);
  nand GNAME1186(G1186,G2345,G7228,G7229);
  nand GNAME1187(G1187,G2345,G7232,G7233);
  nand GNAME1188(G1188,G5216,G5217);
  nand GNAME1189(G1189,G5218,G6772);
  nand GNAME1190(G1190,G1249,G1252,G1253,G1264);
  and GNAME1191(G1191,G1282,G2610);
  nand GNAME1192(G1192,G1773,G1774,G1775,G1776);
  nand GNAME1193(G1193,G4159,G21560);
  not GNAME1194(G1194,G21391);
  and GNAME1195(G1195,G1204,G21391);
  and GNAME1196(G1196,G1197,G1195);
  not GNAME1197(G1197,G21390);
  and GNAME1198(G1198,G1195,G21390);
  not GNAME1199(G1199,G21759);
  and GNAME1200(G1200,G7292,G1194);
  and GNAME1201(G1201,G1197,G21391);
  not GNAME1202(G1202,G35);
  and GNAME1203(G1203,G1201,G2315,G2441);
  not GNAME1204(G1204,G21392);
  or GNAME1205(G1205,G36,G21798);
  not GNAME1206(G1206,G21393);
  not GNAME1207(G1207,G21394);
  not GNAME1208(G1208,G21425);
  not GNAME1209(G1209,G21426);
  not GNAME1210(G1210,G21561);
  not GNAME1211(G1211,G21560);
  not GNAME1212(G1212,G21559);
  not GNAME1213(G1213,G21558);
  nor GNAME1214(G1214,G1212,G1213);
  and GNAME1215(G1215,G21561,G21560);
  and GNAME1216(G1216,G1214,G1215);
  and GNAME1217(G1217,G1210,G21560);
  and GNAME1218(G1218,G1214,G1217);
  and GNAME1219(G1219,G1211,G21561);
  and GNAME1220(G1220,G1214,G1219);
  nor GNAME1221(G1221,G21561,G21560);
  and GNAME1222(G1222,G1214,G1221);
  and GNAME1223(G1223,G1212,G21558);
  nor GNAME1224(G1224,G2348,G2349);
  and GNAME1225(G1225,G1217,G1223);
  and GNAME1226(G1226,G1219,G1223);
  and GNAME1227(G1227,G1221,G1223);
  nor GNAME1228(G1228,G21558,G1212);
  and GNAME1229(G1229,G1215,G1228);
  and GNAME1230(G1230,G1217,G1228);
  and GNAME1231(G1231,G1219,G1228);
  and GNAME1232(G1232,G1221,G1228);
  nor GNAME1233(G1233,G21559,G21558);
  and GNAME1234(G1234,G1215,G1233);
  and GNAME1235(G1235,G1217,G1233);
  and GNAME1236(G1236,G1219,G1233);
  and GNAME1237(G1237,G1221,G1233);
  nand GNAME1238(G1238,G1793,G1794,G1795,G1796);
  nand GNAME1239(G1239,G1797,G1798,G1799,G1800);
  nand GNAME1240(G1240,G1789,G1790,G1791,G1792);
  nor GNAME1241(G1241,G2579,G1240);
  nand GNAME1242(G1242,G1777,G1778,G1779,G1780);
  and GNAME1243(G1243,G1249,G1241);
  nor GNAME1244(G1244,G1238,G1239);
  nand GNAME1245(G1245,G1202,G1276);
  nand GNAME1246(G1246,G1204,G2459);
  nand GNAME1247(G1247,G1243,G1244,G2477,G1248,G2494);
  nand GNAME1248(G1248,G1769,G1770,G1771,G1772);
  nand GNAME1249(G1249,G1781,G1782,G1783,G1784);
  nor GNAME1250(G1250,G1192,G1249);
  and GNAME1251(G1251,G1242,G1239,G1252,G1250);
  nand GNAME1252(G1252,G1785,G1786,G1787,G1788);
  and GNAME1253(G1253,G2494,G2528);
  and GNAME1254(G1254,G1252,G2311,G6746);
  and GNAME1255(G1255,G1202,G2459);
  and GNAME1256(G1256,G2598,G2604,G2605,G1254);
  nand GNAME1257(G1257,G2346,G2606,G2607,G1256);
  nor GNAME1258(G1258,G2596,G1248);
  nor GNAME1259(G1259,G2608,G1239);
  and GNAME1260(G1260,G1249,G2511);
  and GNAME1261(G1261,G1238,G2528);
  and GNAME1262(G1262,G1192,G1248);
  or GNAME1263(G1263,G1523,G1525);
  and GNAME1264(G1264,G2596,G683,G1248);
  nor GNAME1265(G1265,G2477,G1192);
  and GNAME1266(G1266,G1265,G1239,G1241);
  and GNAME1267(G1267,G1266,G1248,G1249);
  nand GNAME1268(G1268,G1801,G8114,G6747,G6748);
  not GNAME1269(G1269,G21428);
  and GNAME1270(G1270,G2597,G21426);
  nand GNAME1271(G1271,G6777,G6778,G2614,G1270);
  not GNAME1272(G1272,G21427);
  and GNAME1273(G1273,G21426,G21427);
  and GNAME1274(G1274,G21428,G1273);
  nor GNAME1275(G1275,G21426,G1269);
  not GNAME1276(G1276,G21797);
  and GNAME1277(G1277,G21427,G21797);
  and GNAME1278(G1278,G1276,G21427);
  nor GNAME1279(G1279,G21426,G2298);
  nor GNAME1280(G1280,G21425,G21427);
  and GNAME1281(G1281,G1209,G1272);
  not GNAME1282(G1282,G7326);
  and GNAME1283(G1283,G1272,G21426);
  not GNAME1284(G1284,G21565);
  not GNAME1285(G1285,G21566);
  not GNAME1286(G1286,G21564);
  not GNAME1287(G1287,G21563);
  and GNAME1288(G1288,G21564,G21565,G21566);
  nor GNAME1289(G1289,G2629,G2637);
  nor GNAME1290(G1290,G21566,G2642);
  and GNAME1291(G1291,G1269,G21425);
  and GNAME1292(G1292,G1269,G21426);
  nor GNAME1293(G1293,G2690,G2298);
  and GNAME1294(G1294,G21563,G1288);
  and GNAME1295(G1295,G1321,G1293);
  and GNAME1296(G1296,G21426,G2511);
  nand GNAME1297(G1297,G1248,G2562);
  or GNAME1298(G1298,G2655,G1544);
  nor GNAME1299(G1299,G21427,G1269);
  not GNAME1300(G1300,G1760);
  nand GNAME1301(G1301,G6783,G6784,G2615,G2649);
  or GNAME1302(G1302,G1526,G2647,G1209,G1269);
  nand GNAME1303(G1303,G2651,G2670);
  nand GNAME1304(G1304,G2633,G2309);
  nand GNAME1305(G1305,G2645,G2643,G2644);
  and GNAME1306(G1306,G1301,G1302);
  nand GNAME1307(G1307,G2667,G2668);
  or GNAME1308(G1308,G1296,G1313);
  nand GNAME1309(G1309,G2640,G2638,G2639);
  nand GNAME1310(G1310,G2249,G2663);
  nand GNAME1311(G1311,G2675,G2676);
  and GNAME1312(G1312,G21426,G2545);
  and GNAME1313(G1313,G2671,G2672);
  nand GNAME1314(G1314,G2664,G2665);
  nand GNAME1315(G1315,G1308,G2684);
  and GNAME1316(G1316,G1739,G2277);
  nor GNAME1317(G1317,G6801,G6807);
  nor GNAME1318(G1318,G2690,G2307);
  nor GNAME1319(G1319,G1310,G6794,G1303);
  and GNAME1320(G1320,G1323,G1321);
  nand GNAME1321(G1321,G1289,G1290);
  nor GNAME1322(G1322,G2286,G1321);
  nand GNAME1323(G1323,G6804,G1319);
  nor GNAME1324(G1324,G1326,G7291);
  and GNAME1325(G1325,G1318,G1);
  and GNAME1326(G1326,G1316,G1317);
  and GNAME1327(G1327,G1531,G2700);
  and GNAME1328(G1328,G1531,G25);
  and GNAME1329(G1329,G1318,G2);
  and GNAME1330(G1330,G1531,G2713);
  and GNAME1331(G1331,G1531,G26);
  and GNAME1332(G1332,G1318,G3);
  and GNAME1333(G1333,G1531,G2726);
  and GNAME1334(G1334,G1531,G27);
  and GNAME1335(G1335,G1318,G4);
  and GNAME1336(G1336,G1531,G2739);
  and GNAME1337(G1337,G1531,G28);
  and GNAME1338(G1338,G1318,G5);
  and GNAME1339(G1339,G1531,G2752);
  and GNAME1340(G1340,G1531,G29);
  and GNAME1341(G1341,G1318,G6);
  and GNAME1342(G1342,G1531,G2765);
  and GNAME1343(G1343,G1531,G30);
  and GNAME1344(G1344,G1318,G7);
  and GNAME1345(G1345,G1531,G2778);
  and GNAME1346(G1346,G1531,G31);
  and GNAME1347(G1347,G1318,G8);
  and GNAME1348(G1348,G1531,G2791);
  and GNAME1349(G1349,G1531,G32);
  nor GNAME1350(G1350,G2642,G1285);
  and GNAME1351(G1351,G1285,G21565);
  and GNAME1352(G1352,G21564,G1351);
  nand GNAME1353(G1353,G21563,G1352);
  and GNAME1354(G1354,G1358,G1293);
  and GNAME1355(G1355,G1315,G1739);
  nor GNAME1356(G1356,G1310,G2258,G6794);
  and GNAME1357(G1357,G1360,G1358);
  nand GNAME1358(G1358,G1289,G1350);
  nor GNAME1359(G1359,G2285,G1358);
  nand GNAME1360(G1360,G6804,G1356);
  nor GNAME1361(G1361,G1362,G7291);
  and GNAME1362(G1362,G1317,G1355);
  or GNAME1363(G1363,G1351,G1365);
  nor GNAME1364(G1364,G21566,G1363);
  and GNAME1365(G1365,G1284,G21566);
  and GNAME1366(G1366,G21564,G1365);
  nand GNAME1367(G1367,G21563,G1366);
  and GNAME1368(G1368,G1372,G1293);
  nor GNAME1369(G1369,G6807,G1728);
  nor GNAME1370(G1370,G1727,G1303,G1310);
  and GNAME1371(G1371,G1374,G1372);
  nand GNAME1372(G1372,G1289,G1364);
  nor GNAME1373(G1373,G2284,G1372);
  nand GNAME1374(G1374,G6804,G1370);
  nor GNAME1375(G1375,G1376,G7291);
  and GNAME1376(G1376,G1316,G1369);
  nor GNAME1377(G1377,G1285,G1363);
  nor GNAME1378(G1378,G1286,G21566,G21565);
  nand GNAME1379(G1379,G21563,G1378);
  and GNAME1380(G1380,G1383,G1293);
  nor GNAME1381(G1381,G1727,G2258,G1310);
  and GNAME1382(G1382,G1385,G1383);
  nand GNAME1383(G1383,G1289,G1377);
  nor GNAME1384(G1384,G2283,G1383);
  nand GNAME1385(G1385,G6804,G1381);
  nor GNAME1386(G1386,G1387,G7291);
  and GNAME1387(G1387,G1355,G1369);
  or GNAME1388(G1388,G2636,G1390);
  nor GNAME1389(G1389,G2629,G1388);
  and GNAME1390(G1390,G21566,G1286,G21565);
  nand GNAME1391(G1391,G21563,G1390);
  and GNAME1392(G1392,G1396,G1293);
  nor GNAME1393(G1393,G1739,G1315);
  nor GNAME1394(G1394,G1303,G2259,G6794);
  and GNAME1395(G1395,G1398,G1396);
  nand GNAME1396(G1396,G1290,G1389);
  nor GNAME1397(G1397,G2282,G1396);
  nand GNAME1398(G1398,G6804,G1394);
  nor GNAME1399(G1399,G1400,G7291);
  and GNAME1400(G1400,G1317,G1393);
  and GNAME1401(G1401,G1286,G1351);
  nand GNAME1402(G1402,G21563,G1401);
  and GNAME1403(G1403,G1407,G1293);
  nor GNAME1404(G1404,G2277,G1739);
  nor GNAME1405(G1405,G6794,G2258,G2259);
  and GNAME1406(G1406,G1409,G1407);
  nand GNAME1407(G1407,G1350,G1389);
  nor GNAME1408(G1408,G2281,G1407);
  nand GNAME1409(G1409,G6804,G1405);
  nor GNAME1410(G1410,G1411,G7291);
  and GNAME1411(G1411,G1317,G1404);
  and GNAME1412(G1412,G1286,G1365);
  nand GNAME1413(G1413,G21563,G1412);
  and GNAME1414(G1414,G1417,G1293);
  nor GNAME1415(G1415,G1727,G2259,G1303);
  and GNAME1416(G1416,G1419,G1417);
  nand GNAME1417(G1417,G1364,G1389);
  nor GNAME1418(G1418,G2280,G1417);
  nand GNAME1419(G1419,G6804,G1415);
  nor GNAME1420(G1420,G1421,G7291);
  and GNAME1421(G1421,G1369,G1393);
  nor GNAME1422(G1422,G21564,G21565,G21566);
  nand GNAME1423(G1423,G21563,G1422);
  and GNAME1424(G1424,G1427,G1293);
  nor GNAME1425(G1425,G1727,G2258,G2259);
  and GNAME1426(G1426,G1429,G1427);
  nand GNAME1427(G1427,G1377,G1389);
  nor GNAME1428(G1428,G2279,G1427);
  nand GNAME1429(G1429,G6804,G1425);
  nor GNAME1430(G1430,G1431,G7291);
  and GNAME1431(G1431,G1369,G1404);
  nor GNAME1432(G1432,G6801,G1729);
  nand GNAME1433(G1433,G2628,G2268);
  nor GNAME1434(G1434,G2637,G1433);
  and GNAME1435(G1435,G1287,G1288);
  and GNAME1436(G1436,G1437,G1439);
  nand GNAME1437(G1437,G1290,G1434);
  nor GNAME1438(G1438,G2276,G1437);
  nand GNAME1439(G1439,G1726,G1319);
  nor GNAME1440(G1440,G1442,G7291);
  and GNAME1441(G1441,G1437,G1293);
  and GNAME1442(G1442,G1316,G1432);
  nand GNAME1443(G1443,G1287,G1352);
  and GNAME1444(G1444,G1445,G1447);
  nand GNAME1445(G1445,G1350,G1434);
  nor GNAME1446(G1446,G2275,G1445);
  nand GNAME1447(G1447,G1726,G1356);
  nor GNAME1448(G1448,G1450,G7291);
  and GNAME1449(G1449,G1445,G1293);
  and GNAME1450(G1450,G1355,G1432);
  nor GNAME1451(G1451,G1728,G1729);
  nand GNAME1452(G1452,G1287,G1366);
  and GNAME1453(G1453,G1454,G1456);
  nand GNAME1454(G1454,G1364,G1434);
  nor GNAME1455(G1455,G2274,G1454);
  nand GNAME1456(G1456,G1726,G1370);
  nor GNAME1457(G1457,G1459,G7291);
  and GNAME1458(G1458,G1454,G1293);
  and GNAME1459(G1459,G1316,G1451);
  nand GNAME1460(G1460,G1287,G1378);
  and GNAME1461(G1461,G1462,G1464);
  nand GNAME1462(G1462,G1377,G1434);
  nor GNAME1463(G1463,G2273,G1462);
  nand GNAME1464(G1464,G1726,G1381);
  nor GNAME1465(G1465,G1467,G7291);
  and GNAME1466(G1466,G1462,G1293);
  and GNAME1467(G1467,G1355,G1451);
  nor GNAME1468(G1468,G1388,G1433);
  nand GNAME1469(G1469,G1287,G1390);
  and GNAME1470(G1470,G1471,G1473);
  nand GNAME1471(G1471,G1290,G1468);
  nor GNAME1472(G1472,G2272,G1471);
  nand GNAME1473(G1473,G1726,G1394);
  nor GNAME1474(G1474,G1476,G7291);
  and GNAME1475(G1475,G1471,G1293);
  and GNAME1476(G1476,G1393,G1432);
  nand GNAME1477(G1477,G1287,G1401);
  and GNAME1478(G1478,G1479,G1481);
  nand GNAME1479(G1479,G1350,G1468);
  nor GNAME1480(G1480,G2271,G1479);
  nand GNAME1481(G1481,G1726,G1405);
  nor GNAME1482(G1482,G1484,G7291);
  and GNAME1483(G1483,G1479,G1293);
  and GNAME1484(G1484,G1404,G1432);
  nand GNAME1485(G1485,G1287,G1412);
  and GNAME1486(G1486,G1487,G1489);
  nand GNAME1487(G1487,G1364,G1468);
  nor GNAME1488(G1488,G2270,G1487);
  nand GNAME1489(G1489,G1726,G1415);
  nor GNAME1490(G1490,G1492,G7291);
  and GNAME1491(G1491,G1487,G1293);
  and GNAME1492(G1492,G1393,G1451);
  nand GNAME1493(G1493,G1287,G1422);
  and GNAME1494(G1494,G1495,G1497);
  nand GNAME1495(G1495,G1377,G1468);
  nor GNAME1496(G1496,G2269,G1495);
  nand GNAME1497(G1497,G1726,G1425);
  nor GNAME1498(G1498,G1500,G7291);
  and GNAME1499(G1499,G1495,G1293);
  and GNAME1500(G1500,G1404,G1451);
  and GNAME1501(G1501,G2596,G2511);
  not GNAME1502(G1502,G8101);
  and GNAME1503(G1503,G1251,G1258);
  nand GNAME1504(G1504,G2545,G1503);
  and GNAME1505(G1505,G1932,G1254,G4105,G4125);
  nor GNAME1506(G1506,G1269,G2332);
  nor GNAME1507(G1507,G21426,G1282);
  not GNAME1508(G1508,G7779);
  and GNAME1509(G1509,G2596,G2562);
  nor GNAME1510(G1510,G2311,G1192,G1252);
  nor GNAME1511(G1511,G2528,G2545);
  and GNAME1512(G1512,G1242,G1250,G1258,G1511);
  and GNAME1513(G1513,G1250,G2579,G1244,G1240,G2477);
  nor GNAME1514(G1514,G2311,G2579,G1248);
  nand GNAME1515(G1515,G1514,G2545,G2477);
  nor GNAME1516(G1516,G2494,G1242);
  nand GNAME1517(G1517,G1192,G1239);
  and GNAME1518(G1518,G1239,G2477);
  and GNAME1519(G1519,G4125,G4126);
  and GNAME1520(G1520,G4124,G2347,G4123);
  and GNAME1521(G1521,G4128,G1519,G1520,G7194,G7195);
  and GNAME1522(G1522,G1933,G1521,G7197,G2322);
  and GNAME1523(G1523,G1192,G1241,G1259,G1260);
  and GNAME1524(G1524,G4113,G4115);
  and GNAME1525(G1525,G1242,G1243,G1261,G1262);
  and GNAME1526(G1526,G6787,G21427);
  nand GNAME1527(G1527,G4116,G4146);
  not GNAME1528(G1528,G7482);
  not GNAME1529(G1529,G7809);
  not GNAME1530(G1530,G7467);
  nand GNAME1531(G1531,G2689,G6781,G6782);
  nand GNAME1532(G1532,G2690,G2338,G4184);
  and GNAME1533(G1533,G1532,G1279);
  and GNAME1534(G1534,G1532,G4186);
  nand GNAME1535(G1535,G1208,G1281);
  nor GNAME1536(G1536,G1543,G1209);
  and GNAME1537(G1537,G4212,G1536);
  and GNAME1538(G1538,G4211,G1536);
  and GNAME1539(G1539,G4210,G1536);
  and GNAME1540(G1540,G1523,G1536);
  nor GNAME1541(G1541,G21426,G1543);
  not GNAME1542(G1542,G21758);
  and GNAME1543(G1543,G4209,G2344);
  and GNAME1544(G1544,G21426,G1248,G1249);
  nand GNAME1545(G1545,G1544,G1266,G1299);
  nor GNAME1546(G1546,G1550,G1722);
  nor GNAME1547(G1547,G1550,G2317);
  nor GNAME1548(G1548,G1550,G2298);
  nor GNAME1549(G1549,G1550,G1269);
  and GNAME1550(G1550,G4405,G5194);
  or GNAME1551(G1551,G1190,G1269);
  nand GNAME1552(G1552,G2297,G1202,G8101);
  nor GNAME1553(G1553,G1555,G1238);
  nor GNAME1554(G1554,G2545,G1555);
  and GNAME1555(G1555,G4567,G4568);
  nand GNAME1556(G1556,G1238,G1503);
  or GNAME1557(G1557,G1269,G1556);
  nand GNAME1558(G1558,G21428,G2459,G2320);
  nor GNAME1559(G1559,G21428,G1561);
  nor GNAME1560(G1560,G1561,G1269);
  and GNAME1561(G1561,G4650,G4651);
  and GNAME1562(G1562,G1248,G1560);
  nand GNAME1563(G1563,G2545,G2511,G1510,G1518);
  and GNAME1564(G1564,G21428,G2325);
  nand GNAME1565(G1565,G4748,G1283);
  nor GNAME1566(G1566,G1501,G1565);
  and GNAME1567(G1567,G1260,G2328);
  nor GNAME1568(G1568,G2311,G1565);
  nor GNAME1569(G1569,G2511,G1565);
  nor GNAME1570(G1570,G2596,G1565);
  and GNAME1571(G1571,G21428,G1525);
  nand GNAME1572(G1572,G683,G1248,G1239,G1510);
  nand GNAME1573(G1573,G4892,G1283);
  nor GNAME1574(G1574,G2562,G1573);
  nor GNAME1575(G1575,G1249,G1573);
  and GNAME1576(G1576,G4990,G4991);
  and GNAME1577(G1577,G1244,G1583,G21426);
  and GNAME1578(G1578,G2460,G1577);
  and GNAME1579(G1579,G1245,G1583,G21426,G1261);
  and GNAME1580(G1580,G4993,G4994);
  and GNAME1581(G1581,G1583,G4996);
  and GNAME1582(G1582,G1583,G1275);
  nand GNAME1583(G1583,G2342,G2343,G2344,G1576);
  and GNAME1584(G1584,G1578,G1276,G1255);
  nor GNAME1585(G1585,G4992,G1580);
  nand GNAME1586(G1586,G2003,G2005,G2007,G2009);
  nand GNAME1587(G1587,G21759,G2330);
  and GNAME1588(G1588,G4988,G4989);
  and GNAME1589(G1589,G1204,G1197);
  nor GNAME1590(G1590,G7776,G7809);
  nor GNAME1591(G1591,G7779,G7824);
  and GNAME1592(G1592,G1590,G1591);
  nor GNAME1593(G1593,G7776,G1529);
  and GNAME1594(G1594,G1591,G1593);
  and GNAME1595(G1595,G1508,G7824);
  and GNAME1596(G1596,G1590,G1595);
  and GNAME1597(G1597,G1593,G1595);
  and GNAME1598(G1598,G1529,G7776);
  and GNAME1599(G1599,G1591,G1598);
  and GNAME1600(G1600,G7776,G7809);
  and GNAME1601(G1601,G1591,G1600);
  and GNAME1602(G1602,G1595,G1598);
  and GNAME1603(G1603,G1595,G1600);
  and GNAME1604(G1604,G7779,G7824);
  and GNAME1605(G1605,G1600,G1604);
  and GNAME1606(G1606,G1598,G1604);
  nor GNAME1607(G1607,G7824,G1508);
  and GNAME1608(G1608,G1600,G1607);
  and GNAME1609(G1609,G1598,G1607);
  and GNAME1610(G1610,G1593,G1604);
  and GNAME1611(G1611,G1590,G1604);
  and GNAME1612(G1612,G1593,G1607);
  and GNAME1613(G1613,G1590,G1607);
  and GNAME1614(G1614,G1624,G1731);
  and GNAME1615(G1615,G1219,G1614);
  and GNAME1616(G1616,G1221,G1614);
  and GNAME1617(G1617,G1215,G1614);
  and GNAME1618(G1618,G1217,G1614);
  and GNAME1619(G1619,G1624,G7244);
  and GNAME1620(G1620,G1219,G1619);
  and GNAME1621(G1621,G1221,G1619);
  and GNAME1622(G1622,G1215,G1619);
  and GNAME1623(G1623,G1217,G1619);
  nand GNAME1624(G1624,G2349,G7240,G7241);
  nor GNAME1625(G1625,G1731,G1624);
  and GNAME1626(G1626,G1217,G1625);
  and GNAME1627(G1627,G1215,G1625);
  and GNAME1628(G1628,G1221,G1625);
  and GNAME1629(G1629,G1219,G1625);
  nor GNAME1630(G1630,G7244,G1624);
  and GNAME1631(G1631,G1217,G1630);
  and GNAME1632(G1632,G1215,G1630);
  and GNAME1633(G1633,G1221,G1630);
  and GNAME1634(G1634,G1219,G1630);
  nor GNAME1635(G1635,G1524,G1193);
  and GNAME1636(G1636,G21561,G1730);
  and GNAME1637(G1637,G1635,G1636);
  and GNAME1638(G1638,G1210,G1730);
  and GNAME1639(G1639,G1635,G1638);
  nor GNAME1640(G1640,G1524,G4160);
  and GNAME1641(G1641,G1636,G1640);
  and GNAME1642(G1642,G1638,G1640);
  nor GNAME1643(G1643,G1730,G1210);
  and GNAME1644(G1644,G1635,G1643);
  nor GNAME1645(G1645,G1730,G21561);
  and GNAME1646(G1646,G1635,G1645);
  and GNAME1647(G1647,G1640,G1643);
  and GNAME1648(G1648,G1640,G1645);
  and GNAME1649(G1649,G1193,G1524);
  and GNAME1650(G1650,G1645,G1649);
  and GNAME1651(G1651,G1643,G1649);
  and GNAME1652(G1652,G4160,G1524);
  and GNAME1653(G1653,G1645,G1652);
  and GNAME1654(G1654,G1643,G1652);
  and GNAME1655(G1655,G1638,G1649);
  and GNAME1656(G1656,G1636,G1649);
  and GNAME1657(G1657,G1638,G1652);
  and GNAME1658(G1658,G1636,G1652);
  nand GNAME1659(G1659,G2477,G2459,G1248);
  nor GNAME1660(G1660,G1238,G1659);
  and GNAME1661(G1661,G1265,G1282,G1238);
  and GNAME1662(G1662,G682,G1248);
  and GNAME1663(G1663,G7443,G7482);
  and GNAME1664(G1664,G7440,G7467);
  and GNAME1665(G1665,G1663,G1664);
  and GNAME1666(G1666,G1530,G7440);
  and GNAME1667(G1667,G1663,G1666);
  and GNAME1668(G1668,G1528,G7443);
  and GNAME1669(G1669,G1664,G1668);
  and GNAME1670(G1670,G1666,G1668);
  nor GNAME1671(G1671,G7440,G1530);
  and GNAME1672(G1672,G1663,G1671);
  nor GNAME1673(G1673,G7467,G7440);
  and GNAME1674(G1674,G1663,G1673);
  and GNAME1675(G1675,G1668,G1671);
  and GNAME1676(G1676,G1668,G1673);
  nor GNAME1677(G1677,G7443,G1528);
  and GNAME1678(G1678,G1664,G1677);
  and GNAME1679(G1679,G1666,G1677);
  nor GNAME1680(G1680,G7482,G7443);
  and GNAME1681(G1681,G1664,G1680);
  and GNAME1682(G1682,G1666,G1680);
  and GNAME1683(G1683,G1671,G1677);
  and GNAME1684(G1684,G1673,G1677);
  and GNAME1685(G1685,G1671,G1680);
  and GNAME1686(G1686,G1673,G1680);
  and GNAME1687(G1687,G7326,G1238,G1265);
  or GNAME1688(G1688,G1217,G1219);
  nor GNAME1689(G1689,G7204,G1688);
  nor GNAME1690(G1690,G2260,G1210);
  and GNAME1691(G1691,G1689,G1690);
  nor GNAME1692(G1692,G21561,G2260);
  and GNAME1693(G1693,G1689,G1692);
  nor GNAME1694(G1694,G4158,G7204);
  and GNAME1695(G1695,G1690,G1694);
  and GNAME1696(G1696,G1692,G1694);
  nor GNAME1697(G1697,G1210,G1527);
  and GNAME1698(G1698,G1689,G1697);
  nor GNAME1699(G1699,G21561,G1527);
  and GNAME1700(G1700,G1689,G1699);
  and GNAME1701(G1701,G1694,G1697);
  and GNAME1702(G1702,G1694,G1699);
  nor GNAME1703(G1703,G1741,G1688);
  and GNAME1704(G1704,G1690,G1703);
  and GNAME1705(G1705,G1692,G1703);
  nor GNAME1706(G1706,G4158,G1741);
  and GNAME1707(G1707,G1690,G1706);
  and GNAME1708(G1708,G1692,G1706);
  and GNAME1709(G1709,G1697,G1703);
  and GNAME1710(G1710,G1699,G1703);
  and GNAME1711(G1711,G1697,G1706);
  and GNAME1712(G1712,G1699,G1706);
  nand GNAME1713(G1713,G21428,G1523);
  nand GNAME1714(G1714,G7326,G1267,G21428);
  and GNAME1715(G1715,G6355,G2303);
  and GNAME1716(G1716,G1297,G6358,G6359,G1519);
  nand GNAME1717(G1717,G2579,G1512);
  nand GNAME1718(G1718,G21428,G1513);
  and GNAME1719(G1719,G6374,G1558);
  nand GNAME1720(G1720,G21428,G1282,G1267);
  and GNAME1721(G1721,G6415,G2303);
  and GNAME1722(G1722,G2307,G2306);
  or GNAME1723(G1723,G1269,G1563);
  nand GNAME1724(G1724,G1280,G1239,G1249);
  nor GNAME1725(G1725,G2296,G21425);
  nand GNAME1726(G1726,G6802,G6803);
  nand GNAME1727(G1727,G6792,G6793);
  nand GNAME1728(G1728,G6799,G6800);
  nand GNAME1729(G1729,G6805,G6806);
  and GNAME1730(G1730,G7210,G7211);
  nand GNAME1731(G1731,G7242,G7243);
  nand GNAME1732(G1732,G6753,G6754);
  nand GNAME1733(G1733,G6755,G6756);
  nand GNAME1734(G1734,G6757,G6758);
  nand GNAME1735(G1735,G6759,G6760);
  nand GNAME1736(G1736,G6770,G6771);
  nand GNAME1737(G1737,G6773,G6774);
  nand GNAME1738(G1738,G6775,G6776);
  and GNAME1739(G1739,G6795,G6796);
  nand GNAME1740(G1740,G7192,G7193);
  nand GNAME1741(G1741,G7202,G7203);
  nand GNAME1742(G1742,G7205,G7206);
  nand GNAME1743(G1743,G7212,G7213);
  nand GNAME1744(G1744,G7214,G7215);
  nand GNAME1745(G1745,G7216,G7217);
  nand GNAME1746(G1746,G7218,G7219);
  nand GNAME1747(G1747,G7226,G7227);
  nand GNAME1748(G1748,G7230,G7231);
  nand GNAME1749(G1749,G7234,G7235);
  nand GNAME1750(G1750,G7236,G7237);
  nand GNAME1751(G1751,G7238,G7239);
  nand GNAME1752(G1752,G7245,G7246);
  nand GNAME1753(G1753,G7247,G7248);
  nand GNAME1754(G1754,G7249,G7250);
  nand GNAME1755(G1755,G7251,G7252);
  nand GNAME1756(G1756,G7253,G7254);
  nand GNAME1757(G1757,G7255,G7256);
  nand GNAME1758(G1758,G7257,G7258);
  nand GNAME1759(G1759,G7259,G7260);
  nand GNAME1760(G1760,G7261,G7262);
  nand GNAME1761(G1761,G7263,G7264);
  nand GNAME1762(G1762,G7265,G7266);
  nand GNAME1763(G1763,G7267,G7268);
  nand GNAME1764(G1764,G7269,G7270);
  nand GNAME1765(G1765,G7271,G7272);
  nand GNAME1766(G1766,G7273,G7274);
  nand GNAME1767(G1767,G7275,G7276);
  nand GNAME1768(G1768,G7277,G7278);
  and GNAME1769(G1769,G2495,G2496,G2497,G2498);
  and GNAME1770(G1770,G2499,G2500,G2501,G2502);
  and GNAME1771(G1771,G2503,G2504,G2505,G2506);
  and GNAME1772(G1772,G2507,G2508,G2509,G2510);
  and GNAME1773(G1773,G2478,G2479,G2480,G2481);
  and GNAME1774(G1774,G2482,G2483,G2484,G2485);
  and GNAME1775(G1775,G2486,G2487,G2488,G2489);
  and GNAME1776(G1776,G2490,G2491,G2492,G2493);
  and GNAME1777(G1777,G2461,G2462,G2463,G2464);
  and GNAME1778(G1778,G2465,G2466,G2467,G2468);
  and GNAME1779(G1779,G2469,G2470,G2471,G2472);
  and GNAME1780(G1780,G2473,G2474,G2475,G2476);
  and GNAME1781(G1781,G2546,G2547,G2548,G2549);
  and GNAME1782(G1782,G2550,G2551,G2552,G2553);
  and GNAME1783(G1783,G2554,G2555,G2556,G2557);
  and GNAME1784(G1784,G2558,G2559,G2560,G2561);
  and GNAME1785(G1785,G2563,G2564,G2565,G2566);
  and GNAME1786(G1786,G2567,G2568,G2569,G2570);
  and GNAME1787(G1787,G2571,G2572,G2573,G2574);
  and GNAME1788(G1788,G2575,G2576,G2577,G2578);
  and GNAME1789(G1789,G2580,G2581,G2582,G2583);
  and GNAME1790(G1790,G2584,G2585,G2586,G2587);
  and GNAME1791(G1791,G2588,G2589,G2590,G2591);
  and GNAME1792(G1792,G2592,G2593,G2594,G2595);
  and GNAME1793(G1793,G2529,G2530,G2531,G2532);
  and GNAME1794(G1794,G2533,G2534,G2535,G2536);
  and GNAME1795(G1795,G2537,G2538,G2539,G2540);
  and GNAME1796(G1796,G2541,G2542,G2543,G2544);
  and GNAME1797(G1797,G2512,G2513,G2514,G2515);
  and GNAME1798(G1798,G2516,G2517,G2518,G2519);
  and GNAME1799(G1799,G2520,G2521,G2522,G2523);
  and GNAME1800(G1800,G2524,G2525,G2526,G2527);
  nor GNAME1801(G1801,G1267,G8112,G1191);
  and GNAME1802(G1802,G6790,G6791);
  and GNAME1803(G1803,G6797,G6798);
  and GNAME1804(G1804,G2706,G2704,G2705);
  and GNAME1805(G1805,G2719,G2717,G2718);
  and GNAME1806(G1806,G2732,G2730,G2731);
  and GNAME1807(G1807,G2745,G2743,G2744);
  and GNAME1808(G1808,G2758,G2756,G2757);
  and GNAME1809(G1809,G2771,G2769,G2770);
  and GNAME1810(G1810,G2784,G2782,G2783);
  and GNAME1811(G1811,G2797,G2795,G2796);
  and GNAME1812(G1812,G2814,G2812,G2813);
  and GNAME1813(G1813,G2824,G2822,G2823);
  and GNAME1814(G1814,G2834,G2832,G2833);
  and GNAME1815(G1815,G2844,G2842,G2843);
  and GNAME1816(G1816,G2854,G2852,G2853);
  and GNAME1817(G1817,G2864,G2862,G2863);
  and GNAME1818(G1818,G2874,G2872,G2873);
  and GNAME1819(G1819,G2884,G2882,G2883);
  and GNAME1820(G1820,G2901,G2899,G2900);
  and GNAME1821(G1821,G2911,G2909,G2910);
  and GNAME1822(G1822,G2921,G2919,G2920);
  and GNAME1823(G1823,G2931,G2929,G2930);
  and GNAME1824(G1824,G2941,G2939,G2940);
  and GNAME1825(G1825,G2951,G2949,G2950);
  and GNAME1826(G1826,G2961,G2959,G2960);
  and GNAME1827(G1827,G2971,G2969,G2970);
  and GNAME1828(G1828,G2988,G2986,G2987);
  and GNAME1829(G1829,G2998,G2996,G2997);
  and GNAME1830(G1830,G3008,G3006,G3007);
  and GNAME1831(G1831,G3018,G3016,G3017);
  and GNAME1832(G1832,G3028,G3026,G3027);
  and GNAME1833(G1833,G3038,G3036,G3037);
  and GNAME1834(G1834,G3048,G3046,G3047);
  and GNAME1835(G1835,G3058,G3056,G3057);
  and GNAME1836(G1836,G3075,G3073,G3074);
  and GNAME1837(G1837,G3085,G3083,G3084);
  and GNAME1838(G1838,G3095,G3093,G3094);
  and GNAME1839(G1839,G3105,G3103,G3104);
  and GNAME1840(G1840,G3115,G3113,G3114);
  and GNAME1841(G1841,G3125,G3123,G3124);
  and GNAME1842(G1842,G3135,G3133,G3134);
  and GNAME1843(G1843,G3145,G3143,G3144);
  and GNAME1844(G1844,G3162,G3160,G3161);
  and GNAME1845(G1845,G3172,G3170,G3171);
  and GNAME1846(G1846,G3182,G3180,G3181);
  and GNAME1847(G1847,G3192,G3190,G3191);
  and GNAME1848(G1848,G3202,G3200,G3201);
  and GNAME1849(G1849,G3212,G3210,G3211);
  and GNAME1850(G1850,G3222,G3220,G3221);
  and GNAME1851(G1851,G3232,G3230,G3231);
  and GNAME1852(G1852,G3249,G3247,G3248);
  and GNAME1853(G1853,G3259,G3257,G3258);
  and GNAME1854(G1854,G3269,G3267,G3268);
  and GNAME1855(G1855,G3279,G3277,G3278);
  and GNAME1856(G1856,G3289,G3287,G3288);
  and GNAME1857(G1857,G3299,G3297,G3298);
  and GNAME1858(G1858,G3309,G3307,G3308);
  and GNAME1859(G1859,G3319,G3317,G3318);
  and GNAME1860(G1860,G3336,G3334,G3335);
  and GNAME1861(G1861,G3346,G3344,G3345);
  and GNAME1862(G1862,G3356,G3354,G3355);
  and GNAME1863(G1863,G3366,G3364,G3365);
  and GNAME1864(G1864,G3376,G3374,G3375);
  and GNAME1865(G1865,G3386,G3384,G3385);
  and GNAME1866(G1866,G3396,G3394,G3395);
  and GNAME1867(G1867,G3406,G3404,G3405);
  and GNAME1868(G1868,G3423,G3421,G3422);
  and GNAME1869(G1869,G3433,G3431,G3432);
  and GNAME1870(G1870,G3443,G3441,G3442);
  and GNAME1871(G1871,G3453,G3451,G3452);
  and GNAME1872(G1872,G3463,G3461,G3462);
  and GNAME1873(G1873,G3473,G3471,G3472);
  and GNAME1874(G1874,G3483,G3481,G3482);
  and GNAME1875(G1875,G3493,G3491,G3492);
  and GNAME1876(G1876,G3510,G3508,G3509);
  and GNAME1877(G1877,G3520,G3518,G3519);
  and GNAME1878(G1878,G3530,G3528,G3529);
  and GNAME1879(G1879,G3540,G3538,G3539);
  and GNAME1880(G1880,G3550,G3548,G3549);
  and GNAME1881(G1881,G3560,G3558,G3559);
  and GNAME1882(G1882,G3570,G3568,G3569);
  and GNAME1883(G1883,G3580,G3578,G3579);
  and GNAME1884(G1884,G3597,G3595,G3596);
  and GNAME1885(G1885,G3607,G3605,G3606);
  and GNAME1886(G1886,G3617,G3615,G3616);
  and GNAME1887(G1887,G3627,G3625,G3626);
  and GNAME1888(G1888,G3637,G3635,G3636);
  and GNAME1889(G1889,G3647,G3645,G3646);
  and GNAME1890(G1890,G3657,G3655,G3656);
  and GNAME1891(G1891,G3667,G3665,G3666);
  and GNAME1892(G1892,G3684,G3682,G3683);
  and GNAME1893(G1893,G3694,G3692,G3693);
  and GNAME1894(G1894,G3704,G3702,G3703);
  and GNAME1895(G1895,G3714,G3712,G3713);
  and GNAME1896(G1896,G3724,G3722,G3723);
  and GNAME1897(G1897,G3734,G3732,G3733);
  and GNAME1898(G1898,G3744,G3742,G3743);
  and GNAME1899(G1899,G3754,G3752,G3753);
  and GNAME1900(G1900,G3771,G3769,G3770);
  and GNAME1901(G1901,G3781,G3779,G3780);
  and GNAME1902(G1902,G3791,G3789,G3790);
  and GNAME1903(G1903,G3801,G3799,G3800);
  and GNAME1904(G1904,G3811,G3809,G3810);
  and GNAME1905(G1905,G3821,G3819,G3820);
  and GNAME1906(G1906,G3831,G3829,G3830);
  and GNAME1907(G1907,G3841,G3839,G3840);
  and GNAME1908(G1908,G3858,G3856,G3857);
  and GNAME1909(G1909,G3868,G3866,G3867);
  and GNAME1910(G1910,G3878,G3876,G3877);
  and GNAME1911(G1911,G3888,G3886,G3887);
  and GNAME1912(G1912,G3898,G3896,G3897);
  and GNAME1913(G1913,G3908,G3906,G3907);
  and GNAME1914(G1914,G3918,G3916,G3917);
  and GNAME1915(G1915,G3928,G3926,G3927);
  and GNAME1916(G1916,G3945,G3943,G3944);
  and GNAME1917(G1917,G3955,G3953,G3954);
  and GNAME1918(G1918,G3965,G3963,G3964);
  and GNAME1919(G1919,G3975,G3973,G3974);
  and GNAME1920(G1920,G3985,G3983,G3984);
  and GNAME1921(G1921,G3995,G3993,G3994);
  and GNAME1922(G1922,G4005,G4003,G4004);
  and GNAME1923(G1923,G4015,G4013,G4014);
  and GNAME1924(G1924,G4032,G4030,G4031);
  and GNAME1925(G1925,G4042,G4040,G4041);
  and GNAME1926(G1926,G4052,G4050,G4051);
  and GNAME1927(G1927,G4062,G4060,G4061);
  and GNAME1928(G1928,G4072,G4070,G4071);
  and GNAME1929(G1929,G4082,G4080,G4081);
  and GNAME1930(G1930,G4092,G4090,G4091);
  and GNAME1931(G1931,G4102,G4100,G4101);
  and GNAME1932(G1932,G4103,G2347,G1517);
  and GNAME1933(G1933,G7196,G1247,G7200,G7201);
  and GNAME1934(G1934,G4141,G4137,G4140);
  and GNAME1935(G1935,G4152,G4148,G4151);
  and GNAME1936(G1936,G4167,G4165,G4162);
  and GNAME1937(G1937,G2323,G2324);
  and GNAME1938(G1938,G4215,G4218,G4214);
  and GNAME1939(G1939,G4221,G4224,G4220);
  and GNAME1940(G1940,G4227,G4230,G4226);
  and GNAME1941(G1941,G4233,G4236,G4232);
  and GNAME1942(G1942,G4239,G4242,G4238);
  and GNAME1943(G1943,G4245,G4248,G4244);
  and GNAME1944(G1944,G4251,G4254,G4250);
  and GNAME1945(G1945,G4257,G4260,G4256);
  and GNAME1946(G1946,G4263,G4266,G4262);
  and GNAME1947(G1947,G4269,G4272,G4268);
  and GNAME1948(G1948,G4275,G4278,G4274);
  and GNAME1949(G1949,G4281,G4284,G4280);
  and GNAME1950(G1950,G4287,G4290,G4286);
  and GNAME1951(G1951,G4293,G4296,G4292);
  and GNAME1952(G1952,G4299,G4302,G4298);
  and GNAME1953(G1953,G4305,G4308,G4304);
  and GNAME1954(G1954,G4311,G4314,G4310);
  and GNAME1955(G1955,G4317,G4320,G4316);
  and GNAME1956(G1956,G4323,G4326,G4322);
  and GNAME1957(G1957,G4329,G4332,G4328);
  and GNAME1958(G1958,G4335,G4338,G4334);
  and GNAME1959(G1959,G4341,G4344,G4340);
  and GNAME1960(G1960,G4347,G4350,G4346);
  and GNAME1961(G1961,G4353,G4356,G4352);
  and GNAME1962(G1962,G4359,G4362,G4358);
  and GNAME1963(G1963,G4365,G4368,G4364);
  and GNAME1964(G1964,G4371,G4374,G4370);
  and GNAME1965(G1965,G4377,G4380,G4376);
  and GNAME1966(G1966,G4383,G4386,G4382);
  and GNAME1967(G1967,G4389,G4392,G4388);
  and GNAME1968(G1968,G4395,G4398,G4394);
  and GNAME1969(G1969,G4401,G4404,G4400);
  and GNAME1970(G1970,G5003,G5000,G5002);
  and GNAME1971(G1971,G5009,G5006,G5008);
  and GNAME1972(G1972,G5015,G5012,G5014);
  and GNAME1973(G1973,G5021,G5018,G5020);
  and GNAME1974(G1974,G5027,G2333,G5026);
  and GNAME1975(G1975,G5033,G2333,G5032);
  and GNAME1976(G1976,G5039,G2333,G5038);
  and GNAME1977(G1977,G5045,G2333,G5044);
  and GNAME1978(G1978,G5051,G2333,G5050);
  and GNAME1979(G1979,G5057,G2333,G5056);
  and GNAME1980(G1980,G5063,G2333,G5062);
  and GNAME1981(G1981,G5069,G2333,G5068);
  and GNAME1982(G1982,G5075,G2333,G5074);
  and GNAME1983(G1983,G5081,G2333,G5080);
  and GNAME1984(G1984,G5087,G2333,G5086);
  and GNAME1985(G1985,G5093,G2333,G5092);
  and GNAME1986(G1986,G5099,G2333,G5098);
  and GNAME1987(G1987,G5105,G2333,G5104);
  and GNAME1988(G1988,G5111,G2333,G5110);
  and GNAME1989(G1989,G5117,G2333,G5116);
  and GNAME1990(G1990,G5123,G5120,G5122);
  and GNAME1991(G1991,G5129,G5126,G5128);
  and GNAME1992(G1992,G5135,G5132,G5134);
  and GNAME1993(G1993,G5141,G5138,G5140);
  and GNAME1994(G1994,G5147,G5144,G5146);
  and GNAME1995(G1995,G5153,G5151,G5152);
  and GNAME1996(G1996,G5159,G5157,G5158);
  and GNAME1997(G1997,G5165,G5163,G5164);
  and GNAME1998(G1998,G5171,G5169,G5170);
  and GNAME1999(G1999,G5177,G5175,G5176);
  and GNAME2000(G2000,G5183,G5181,G5182);
  and GNAME2001(G2001,G5189,G5187,G5188);
  or GNAME2002(G2002,G21398,G21397,G21396,G21395);
  nor GNAME2003(G2003,G2002,G21399,G21400,G21401,G21402);
  or GNAME2004(G2004,G21406,G21405,G21404,G21403);
  nor GNAME2005(G2005,G2004,G21407,G21408,G21409,G21410);
  or GNAME2006(G2006,G21414,G21413,G21412,G21411);
  nor GNAME2007(G2007,G2006,G21415,G21416,G21417,G21418);
  or GNAME2008(G2008,G21422,G21421,G21420,G21419);
  nor GNAME2009(G2009,G2008,G5190,G21423,G21424);
  and GNAME2010(G2010,G5220,G5221,G5222,G5223);
  and GNAME2011(G2011,G5224,G5225,G5226,G5227);
  and GNAME2012(G2012,G5228,G5229,G5230,G5231);
  and GNAME2013(G2013,G5232,G5233,G5234,G5235);
  and GNAME2014(G2014,G5236,G5237,G5238,G5239);
  and GNAME2015(G2015,G5240,G5241,G5242,G5243);
  and GNAME2016(G2016,G5244,G5245,G5246,G5247);
  and GNAME2017(G2017,G5248,G5249,G5250,G5251);
  and GNAME2018(G2018,G5252,G5253,G5254,G5255);
  and GNAME2019(G2019,G5256,G5257,G5258,G5259);
  and GNAME2020(G2020,G5260,G5261,G5262,G5263);
  and GNAME2021(G2021,G5264,G5265,G5266,G5267);
  and GNAME2022(G2022,G5268,G5269,G5270,G5271);
  and GNAME2023(G2023,G5272,G5273,G5274,G5275);
  and GNAME2024(G2024,G5276,G5277,G5278,G5279);
  and GNAME2025(G2025,G5280,G5281,G5282,G5283);
  and GNAME2026(G2026,G5284,G5285,G5286,G5287);
  and GNAME2027(G2027,G5288,G5289,G5290,G5291);
  and GNAME2028(G2028,G5292,G5293,G5294,G5295);
  and GNAME2029(G2029,G5296,G5297,G5298,G5299);
  and GNAME2030(G2030,G5300,G5301,G5302,G5303);
  and GNAME2031(G2031,G5304,G5305,G5306,G5307);
  and GNAME2032(G2032,G5308,G5309,G5310,G5311);
  and GNAME2033(G2033,G5312,G5313,G5314,G5315);
  and GNAME2034(G2034,G5316,G5317,G5318,G5319);
  and GNAME2035(G2035,G5320,G5321,G5322,G5323);
  and GNAME2036(G2036,G5324,G5325,G5326,G5327);
  and GNAME2037(G2037,G5328,G5329,G5330,G5331);
  and GNAME2038(G2038,G5332,G5333,G5334,G5335);
  and GNAME2039(G2039,G5336,G5337,G5338,G5339);
  and GNAME2040(G2040,G5340,G5341,G5342,G5343);
  and GNAME2041(G2041,G5344,G5345,G5346,G5347);
  and GNAME2042(G2042,G5348,G5349,G5350,G5351);
  and GNAME2043(G2043,G5352,G5353,G5354,G5355);
  and GNAME2044(G2044,G5356,G5357,G5358,G5359);
  and GNAME2045(G2045,G5360,G5361,G5362,G5363);
  and GNAME2046(G2046,G5364,G5365,G5366,G5367);
  and GNAME2047(G2047,G5368,G5369,G5370,G5371);
  and GNAME2048(G2048,G5372,G5373,G5374,G5375);
  and GNAME2049(G2049,G5376,G5377,G5378,G5379);
  and GNAME2050(G2050,G5380,G5381,G5382,G5383);
  and GNAME2051(G2051,G5384,G5385,G5386,G5387);
  and GNAME2052(G2052,G5388,G5389,G5390,G5391);
  and GNAME2053(G2053,G5392,G5393,G5394,G5395);
  and GNAME2054(G2054,G5396,G5397,G5398,G5399);
  and GNAME2055(G2055,G5400,G5401,G5402,G5403);
  and GNAME2056(G2056,G5404,G5405,G5406,G5407);
  and GNAME2057(G2057,G5408,G5409,G5410,G5411);
  and GNAME2058(G2058,G5412,G5413,G5414,G5415);
  and GNAME2059(G2059,G5416,G5417,G5418,G5419);
  and GNAME2060(G2060,G5420,G5421,G5422,G5423);
  and GNAME2061(G2061,G5424,G5425,G5426,G5427);
  and GNAME2062(G2062,G5428,G5429,G5430,G5431);
  and GNAME2063(G2063,G5432,G5433,G5434,G5435);
  and GNAME2064(G2064,G5436,G5437,G5438,G5439);
  and GNAME2065(G2065,G5440,G5441,G5442,G5443);
  and GNAME2066(G2066,G5444,G5445,G5446,G5447);
  and GNAME2067(G2067,G5448,G5449,G5450,G5451);
  and GNAME2068(G2068,G5452,G5453,G5454,G5455);
  and GNAME2069(G2069,G5456,G5457,G5458,G5459);
  and GNAME2070(G2070,G5460,G5461,G5462,G5463);
  and GNAME2071(G2071,G5464,G5465,G5466,G5467);
  and GNAME2072(G2072,G5468,G5469,G5470,G5471);
  and GNAME2073(G2073,G5472,G5473,G5474,G5475);
  and GNAME2074(G2074,G5476,G5477,G5478,G5479);
  and GNAME2075(G2075,G5480,G5481,G5482,G5483);
  and GNAME2076(G2076,G5484,G5485,G5486,G5487);
  and GNAME2077(G2077,G5488,G5489,G5490,G5491);
  and GNAME2078(G2078,G5493,G5494,G5495,G5496);
  and GNAME2079(G2079,G5497,G5498,G5499,G5500);
  and GNAME2080(G2080,G5501,G5502,G5503,G5504);
  and GNAME2081(G2081,G5505,G5506,G5507,G5508);
  and GNAME2082(G2082,G5510,G5511,G5512,G5513);
  and GNAME2083(G2083,G5514,G5515,G5516,G5517);
  and GNAME2084(G2084,G5518,G5519,G5520,G5521);
  and GNAME2085(G2085,G5522,G5523,G5524,G5525);
  and GNAME2086(G2086,G5527,G5528,G5529,G5530);
  and GNAME2087(G2087,G5531,G5532,G5533,G5534);
  and GNAME2088(G2088,G5535,G5536,G5537,G5538);
  and GNAME2089(G2089,G5539,G5540,G5541,G5542);
  and GNAME2090(G2090,G5544,G5545,G5546,G5547);
  and GNAME2091(G2091,G5548,G5549,G5550,G5551);
  and GNAME2092(G2092,G5552,G5553,G5554,G5555);
  and GNAME2093(G2093,G5556,G5557,G5558,G5559);
  and GNAME2094(G2094,G5561,G5562,G5563,G5564);
  and GNAME2095(G2095,G5565,G5566,G5567,G5568);
  and GNAME2096(G2096,G5569,G5570,G5571,G5572);
  and GNAME2097(G2097,G5573,G5574,G5575,G5576);
  and GNAME2098(G2098,G5578,G5579,G5580,G5581);
  and GNAME2099(G2099,G5582,G5583,G5584,G5585);
  and GNAME2100(G2100,G5586,G5587,G5588,G5589);
  and GNAME2101(G2101,G5590,G5591,G5592,G5593);
  and GNAME2102(G2102,G5595,G5596,G5597,G5598);
  and GNAME2103(G2103,G5599,G5600,G5601,G5602);
  and GNAME2104(G2104,G5603,G5604,G5605,G5606);
  and GNAME2105(G2105,G5607,G5608,G5609,G5610);
  and GNAME2106(G2106,G5612,G5613,G5614,G5615);
  and GNAME2107(G2107,G5616,G5617,G5618,G5619);
  and GNAME2108(G2108,G5620,G5621,G5622,G5623);
  and GNAME2109(G2109,G5624,G5625,G5626,G5627);
  and GNAME2110(G2110,G5629,G5630,G5631,G5632);
  and GNAME2111(G2111,G5633,G5634,G5635,G5636);
  and GNAME2112(G2112,G5637,G5638,G5639,G5640);
  and GNAME2113(G2113,G5641,G5642,G5643,G5644);
  and GNAME2114(G2114,G5646,G5647,G5648,G5649);
  and GNAME2115(G2115,G5650,G5651,G5652,G5653);
  and GNAME2116(G2116,G5654,G5655,G5656,G5657);
  and GNAME2117(G2117,G5658,G5659,G5660,G5661);
  and GNAME2118(G2118,G5663,G5664,G5665,G5666);
  and GNAME2119(G2119,G5667,G5668,G5669,G5670);
  and GNAME2120(G2120,G5671,G5672,G5673,G5674);
  and GNAME2121(G2121,G5675,G5676,G5677,G5678);
  and GNAME2122(G2122,G5680,G5681,G5682,G5683);
  and GNAME2123(G2123,G5684,G5685,G5686,G5687);
  and GNAME2124(G2124,G5688,G5689,G5690,G5691);
  and GNAME2125(G2125,G5692,G5693,G5694,G5695);
  and GNAME2126(G2126,G5697,G5698,G5699,G5700);
  and GNAME2127(G2127,G5701,G5702,G5703,G5704);
  and GNAME2128(G2128,G5705,G5706,G5707,G5708);
  and GNAME2129(G2129,G5709,G5710,G5711,G5712);
  and GNAME2130(G2130,G5714,G5715,G5716,G5717);
  and GNAME2131(G2131,G5718,G5719,G5720,G5721);
  and GNAME2132(G2132,G5722,G5723,G5724,G5725);
  and GNAME2133(G2133,G5726,G5727,G5728,G5729);
  and GNAME2134(G2134,G5731,G5732,G5733,G5734);
  and GNAME2135(G2135,G5735,G5736,G5737,G5738);
  and GNAME2136(G2136,G5739,G5740,G5741,G5742);
  and GNAME2137(G2137,G5743,G5744,G5745,G5746);
  and GNAME2138(G2138,G2596,G5907,G5908);
  and GNAME2139(G2139,G5926,G5927,G5928,G5929);
  and GNAME2140(G2140,G5930,G5931,G5932,G5933);
  and GNAME2141(G2141,G5934,G5935,G5936,G5937);
  and GNAME2142(G2142,G5938,G5939,G5940,G5941);
  and GNAME2143(G2143,G5943,G5944,G5945,G5946);
  and GNAME2144(G2144,G5947,G5948,G5949,G5950);
  and GNAME2145(G2145,G5951,G5952,G5953,G5954);
  and GNAME2146(G2146,G5955,G5956,G5957,G5958);
  and GNAME2147(G2147,G5909,G5910,G5911,G5912);
  and GNAME2148(G2148,G5913,G5914,G5915,G5916);
  and GNAME2149(G2149,G5917,G5918,G5919,G5920);
  and GNAME2150(G2150,G5921,G5922,G5923,G5924);
  and GNAME2151(G2151,G5981,G5982,G5983,G5984);
  and GNAME2152(G2152,G5985,G5986,G5987,G5988);
  and GNAME2153(G2153,G5989,G5990,G5991,G5992);
  and GNAME2154(G2154,G5993,G5994,G5995,G5996);
  and GNAME2155(G2155,G5998,G5999,G6000,G6001);
  and GNAME2156(G2156,G6002,G6003,G6004,G6005);
  and GNAME2157(G2157,G6006,G6007,G6008,G6009);
  and GNAME2158(G2158,G6010,G6011,G6012,G6013);
  and GNAME2159(G2159,G5964,G5965,G5966,G5967);
  and GNAME2160(G2160,G5968,G5969,G5970,G5971);
  and GNAME2161(G2161,G5972,G5973,G5974,G5975);
  and GNAME2162(G2162,G5976,G5977,G5978,G5979);
  and GNAME2163(G2163,G6036,G6037,G6038,G6039);
  and GNAME2164(G2164,G6040,G6041,G6042,G6043);
  and GNAME2165(G2165,G6044,G6045,G6046,G6047);
  and GNAME2166(G2166,G6048,G6049,G6050,G6051);
  and GNAME2167(G2167,G6053,G6054,G6055,G6056);
  and GNAME2168(G2168,G6057,G6058,G6059,G6060);
  and GNAME2169(G2169,G6061,G6062,G6063,G6064);
  and GNAME2170(G2170,G6065,G6066,G6067,G6068);
  and GNAME2171(G2171,G6019,G6020,G6021,G6022);
  and GNAME2172(G2172,G6023,G6024,G6025,G6026);
  and GNAME2173(G2173,G6027,G6028,G6029,G6030);
  and GNAME2174(G2174,G6031,G6032,G6033,G6034);
  and GNAME2175(G2175,G6091,G6092,G6093,G6094);
  and GNAME2176(G2176,G6095,G6096,G6097,G6098);
  and GNAME2177(G2177,G6099,G6100,G6101,G6102);
  and GNAME2178(G2178,G6103,G6104,G6105,G6106);
  and GNAME2179(G2179,G6108,G6109,G6110,G6111);
  and GNAME2180(G2180,G6112,G6113,G6114,G6115);
  and GNAME2181(G2181,G6116,G6117,G6118,G6119);
  and GNAME2182(G2182,G6120,G6121,G6122,G6123);
  and GNAME2183(G2183,G6074,G6075,G6076,G6077);
  and GNAME2184(G2184,G6078,G6079,G6080,G6081);
  and GNAME2185(G2185,G6082,G6083,G6084,G6085);
  and GNAME2186(G2186,G6086,G6087,G6088,G6089);
  and GNAME2187(G2187,G6147,G6148,G6149,G6150);
  and GNAME2188(G2188,G6151,G6152,G6153,G6154);
  and GNAME2189(G2189,G6155,G6156,G6157,G6158);
  and GNAME2190(G2190,G6159,G6160,G6161,G6162);
  and GNAME2191(G2191,G6164,G6165,G6166,G6167);
  and GNAME2192(G2192,G6168,G6169,G6170,G6171);
  and GNAME2193(G2193,G6172,G6173,G6174,G6175);
  and GNAME2194(G2194,G6176,G6177,G6178,G6179);
  and GNAME2195(G2195,G6130,G6131,G6132,G6133);
  and GNAME2196(G2196,G6134,G6135,G6136,G6137);
  and GNAME2197(G2197,G6138,G6139,G6140,G6141);
  and GNAME2198(G2198,G6142,G6143,G6144,G6145);
  and GNAME2199(G2199,G6203,G6204,G6205,G6206);
  and GNAME2200(G2200,G6207,G6208,G6209,G6210);
  and GNAME2201(G2201,G6211,G6212,G6213,G6214);
  and GNAME2202(G2202,G6215,G6216,G6217,G6218);
  and GNAME2203(G2203,G6220,G6221,G6222,G6223);
  and GNAME2204(G2204,G6224,G6225,G6226,G6227);
  and GNAME2205(G2205,G6228,G6229,G6230,G6231);
  and GNAME2206(G2206,G6232,G6233,G6234,G6235);
  and GNAME2207(G2207,G6186,G6187,G6188,G6189);
  and GNAME2208(G2208,G6190,G6191,G6192,G6193);
  and GNAME2209(G2209,G6194,G6195,G6196,G6197);
  and GNAME2210(G2210,G6198,G6199,G6200,G6201);
  and GNAME2211(G2211,G6241,G2310,G6237);
  and GNAME2212(G2212,G6259,G6260,G6261,G6262);
  and GNAME2213(G2213,G6263,G6264,G6265,G6266);
  and GNAME2214(G2214,G6267,G6268,G6269,G6270);
  and GNAME2215(G2215,G6271,G6272,G6273,G6274);
  and GNAME2216(G2216,G6276,G6277,G6278,G6279);
  and GNAME2217(G2217,G6280,G6281,G6282,G6283);
  and GNAME2218(G2218,G6284,G6285,G6286,G6287);
  and GNAME2219(G2219,G6288,G6289,G6290,G6291);
  and GNAME2220(G2220,G6242,G6243,G6244,G6245);
  and GNAME2221(G2221,G6246,G6247,G6248,G6249);
  and GNAME2222(G2222,G6250,G6251,G6252,G6253);
  and GNAME2223(G2223,G6254,G6255,G6256,G6257);
  and GNAME2224(G2224,G2312,G1659,G6293,G6297);
  and GNAME2225(G2225,G6315,G6316,G6317,G6318);
  and GNAME2226(G2226,G6319,G6320,G6321,G6322);
  and GNAME2227(G2227,G6323,G6324,G6325,G6326);
  and GNAME2228(G2228,G6327,G6328,G6329,G6330);
  and GNAME2229(G2229,G6332,G6333,G6334,G6335);
  and GNAME2230(G2230,G6336,G6337,G6338,G6339);
  and GNAME2231(G2231,G6340,G6341,G6342,G6343);
  and GNAME2232(G2232,G6344,G6345,G6346,G6347);
  and GNAME2233(G2233,G6298,G6299,G6300,G6301);
  and GNAME2234(G2234,G6302,G6303,G6304,G6305);
  and GNAME2235(G2235,G6306,G6307,G6308,G6309);
  and GNAME2236(G2236,G6310,G6311,G6312,G6313);
  and GNAME2237(G2237,G2310,G2311,G6349,G6353);
  and GNAME2238(G2238,G6356,G6357);
  and GNAME2239(G2239,G2253,G1252,G7280,G6361);
  and GNAME2240(G2240,G2319,G2322,G6368,G6369);
  and GNAME2241(G2241,G2305,G2299,G6376);
  and GNAME2242(G2242,G2317,G1723,G1557);
  and GNAME2243(G2243,G6528,G6526,G6527);
  and GNAME2244(G2244,G6576,G6577,G6575,G6573,G6574);
  and GNAME2245(G2245,G6635,G6636,G6634,G6632,G6633);
  and GNAME2246(G2246,G6694,G6695,G6697,G6696,G6692);
  and GNAME2247(G2247,G6703,G6704,G6706,G6705,G6701);
  and GNAME2248(G2248,G2632,G2630,G2631);
  nand GNAME2249(G2249,G2654,G1309,G2653);
  and GNAME2250(G2250,G2660,G2661);
  nand GNAME2251(G2251,G2679,G2680);
  nand GNAME2252(G2252,G4112,G2338,G2350);
  nand GNAME2253(G2253,G1238,G2511);
  and GNAME2254(G2254,G1215,G2511);
  and GNAME2255(G2255,G1576,G5206,G5207);
  and GNAME2256(G2256,G1535,G1576);
  nand GNAME2257(G2257,G1505,G4110,G4111);
  not GNAME2258(G2258,G1303);
  not GNAME2259(G2259,G1310);
  not GNAME2260(G2260,G1527);
  not GNAME2261(G2261,G1493);
  not GNAME2262(G2262,G1485);
  not GNAME2263(G2263,G1477);
  not GNAME2264(G2264,G1469);
  not GNAME2265(G2265,G1460);
  not GNAME2266(G2266,G1452);
  not GNAME2267(G2267,G1443);
  not GNAME2268(G2268,G1435);
  not GNAME2269(G2269,G1497);
  not GNAME2270(G2270,G1489);
  not GNAME2271(G2271,G1481);
  not GNAME2272(G2272,G1473);
  not GNAME2273(G2273,G1464);
  not GNAME2274(G2274,G1456);
  not GNAME2275(G2275,G1447);
  not GNAME2276(G2276,G1439);
  not GNAME2277(G2277,G1315);
  not GNAME2278(G2278,G1288);
  not GNAME2279(G2279,G1429);
  not GNAME2280(G2280,G1419);
  not GNAME2281(G2281,G1409);
  not GNAME2282(G2282,G1398);
  not GNAME2283(G2283,G1385);
  not GNAME2284(G2284,G1374);
  not GNAME2285(G2285,G1360);
  not GNAME2286(G2286,G1323);
  not GNAME2287(G2287,G1423);
  not GNAME2288(G2288,G1413);
  not GNAME2289(G2289,G1402);
  not GNAME2290(G2290,G1391);
  not GNAME2291(G2291,G1379);
  not GNAME2292(G2292,G1367);
  not GNAME2293(G2293,G1353);
  not GNAME2294(G2294,G1294);
  nand GNAME2295(G2295,G1261,G1280);
  not GNAME2296(G2296,G1724);
  not GNAME2297(G2297,G1551);
  not GNAME2298(G2298,G1278);
  or GNAME2299(G2299,G1269,G1572);
  not GNAME2300(G2300,G1713);
  nand GNAME2301(G2301,G1512,G2459,G21428);
  not GNAME2302(G2302,G1723);
  not GNAME2303(G2303,G1564);
  or GNAME2304(G2304,G2545,G1714);
  nand GNAME2305(G2305,G21428,G1662,G1243,G1239,G2494);
  not GNAME2306(G2306,G1292);
  not GNAME2307(G2307,G1277);
  not GNAME2308(G2308,G1557);
  nand GNAME2309(G2309,G683,G1299);
  not GNAME2310(G2310,G1262);
  not GNAME2311(G2311,G1509);
  not GNAME2312(G2312,G683);
  not GNAME2313(G2313,G1195);
  nand GNAME2314(G2314,G1202,G36);
  or GNAME2315(G2315,G35,G788);
  or GNAME2316(G2316,G35,G1205);
  not GNAME2317(G2317,G1281);
  not GNAME2318(G2318,G1525);
  nand GNAME2319(G2319,G1260,G1266);
  not GNAME2320(G2320,G1247);
  nand GNAME2321(G2321,G1248,G1513);
  or GNAME2322(G2322,G1192,G1515);
  nand GNAME2323(G2323,G1516,G1244,G1514);
  nand GNAME2324(G2324,G1514,G1192,G1259);
  not GNAME2325(G2325,G1504);
  nand GNAME2326(G2326,G2511,G1513);
  or GNAME2327(G2327,G1515,G1517);
  not GNAME2328(G2328,G1565);
  not GNAME2329(G2329,G1261);
  not GNAME2330(G2330,G1586);
  or GNAME2331(G2331,G1272,G7442,G4992);
  not GNAME2332(G2332,G1283);
  nand GNAME2333(G2333,G1583,G1272,G1269);
  nand GNAME2334(G2334,G1246,G1577);
  not GNAME2335(G2335,G1198);
  not GNAME2336(G2336,G1196);
  and GNAME2337(G2337,G1312,G1239,G1583);
  nand GNAME2338(G2338,G1274,G21795);
  nand GNAME2339(G2339,G1542,G1206,G1207,G2330);
  not GNAME2340(G2340,G2254);
  nand GNAME2341(G2341,G35,G1275);
  nand GNAME2342(G2342,G1269,G1279);
  nand GNAME2343(G2343,G1281,G21425,G21428);
  or GNAME2344(G2344,G21428,G1535);
  nand GNAME2345(G2345,G1194,G1589);
  nand GNAME2346(G2346,G2545,G1202,G1240);
  nand GNAME2347(G2347,G1242,G1253);
  not GNAME2348(G2348,G1215);
  not GNAME2349(G2349,G1223);
  not GNAME2350(G2350,G1291);
  nand GNAME2351(G2351,G1196,G21789);
  nand GNAME2352(G2352,G1198,G21788);
  nand GNAME2353(G2353,G2313,G21360);
  nand GNAME2354(G2354,G1196,G21788);
  nand GNAME2355(G2355,G1198,G21787);
  nand GNAME2356(G2356,G2313,G21361);
  nand GNAME2357(G2357,G1196,G21787);
  nand GNAME2358(G2358,G1198,G21786);
  nand GNAME2359(G2359,G2313,G21362);
  nand GNAME2360(G2360,G1196,G21786);
  nand GNAME2361(G2361,G1198,G21785);
  nand GNAME2362(G2362,G2313,G21363);
  nand GNAME2363(G2363,G1196,G21785);
  nand GNAME2364(G2364,G1198,G21784);
  nand GNAME2365(G2365,G2313,G21364);
  nand GNAME2366(G2366,G1196,G21784);
  nand GNAME2367(G2367,G1198,G21783);
  nand GNAME2368(G2368,G2313,G21365);
  nand GNAME2369(G2369,G1196,G21783);
  nand GNAME2370(G2370,G1198,G21782);
  nand GNAME2371(G2371,G2313,G21366);
  nand GNAME2372(G2372,G1196,G21782);
  nand GNAME2373(G2373,G1198,G21781);
  nand GNAME2374(G2374,G2313,G21367);
  nand GNAME2375(G2375,G1196,G21781);
  nand GNAME2376(G2376,G1198,G21780);
  nand GNAME2377(G2377,G2313,G21368);
  nand GNAME2378(G2378,G1196,G21780);
  nand GNAME2379(G2379,G1198,G21779);
  nand GNAME2380(G2380,G2313,G21369);
  nand GNAME2381(G2381,G1196,G21779);
  nand GNAME2382(G2382,G1198,G21778);
  nand GNAME2383(G2383,G2313,G21370);
  nand GNAME2384(G2384,G1196,G21778);
  nand GNAME2385(G2385,G1198,G21777);
  nand GNAME2386(G2386,G2313,G21371);
  nand GNAME2387(G2387,G1196,G21777);
  nand GNAME2388(G2388,G1198,G21776);
  nand GNAME2389(G2389,G2313,G21372);
  nand GNAME2390(G2390,G1196,G21776);
  nand GNAME2391(G2391,G1198,G21775);
  nand GNAME2392(G2392,G2313,G21373);
  nand GNAME2393(G2393,G1196,G21775);
  nand GNAME2394(G2394,G1198,G21774);
  nand GNAME2395(G2395,G2313,G21374);
  nand GNAME2396(G2396,G1196,G21774);
  nand GNAME2397(G2397,G1198,G21773);
  nand GNAME2398(G2398,G2313,G21375);
  nand GNAME2399(G2399,G1196,G21773);
  nand GNAME2400(G2400,G1198,G21772);
  nand GNAME2401(G2401,G2313,G21376);
  nand GNAME2402(G2402,G1196,G21772);
  nand GNAME2403(G2403,G1198,G21771);
  nand GNAME2404(G2404,G2313,G21377);
  nand GNAME2405(G2405,G1196,G21771);
  nand GNAME2406(G2406,G1198,G21770);
  nand GNAME2407(G2407,G2313,G21378);
  nand GNAME2408(G2408,G1196,G21770);
  nand GNAME2409(G2409,G1198,G21769);
  nand GNAME2410(G2410,G2313,G21379);
  nand GNAME2411(G2411,G1196,G21769);
  nand GNAME2412(G2412,G1198,G21768);
  nand GNAME2413(G2413,G2313,G21380);
  nand GNAME2414(G2414,G1196,G21768);
  nand GNAME2415(G2415,G1198,G21767);
  nand GNAME2416(G2416,G2313,G21381);
  nand GNAME2417(G2417,G1196,G21767);
  nand GNAME2418(G2418,G1198,G21766);
  nand GNAME2419(G2419,G2313,G21382);
  nand GNAME2420(G2420,G1196,G21766);
  nand GNAME2421(G2421,G1198,G21765);
  nand GNAME2422(G2422,G2313,G21383);
  nand GNAME2423(G2423,G1196,G21765);
  nand GNAME2424(G2424,G1198,G21764);
  nand GNAME2425(G2425,G2313,G21384);
  nand GNAME2426(G2426,G1196,G21764);
  nand GNAME2427(G2427,G1198,G21763);
  nand GNAME2428(G2428,G2313,G21385);
  nand GNAME2429(G2429,G1196,G21763);
  nand GNAME2430(G2430,G1198,G21762);
  nand GNAME2431(G2431,G2313,G21386);
  nand GNAME2432(G2432,G1196,G21762);
  nand GNAME2433(G2433,G1198,G21761);
  nand GNAME2434(G2434,G2313,G21387);
  nand GNAME2435(G2435,G1196,G21761);
  nand GNAME2436(G2436,G1198,G21760);
  nand GNAME2437(G2437,G2313,G21388);
  nand GNAME2438(G2438,G1196,G21760);
  nand GNAME2439(G2439,G1198,G21759);
  nand GNAME2440(G2440,G2313,G21389);
  nand GNAME2441(G2441,G35,G33,G1201);
  nand GNAME2442(G2442,G6743,G6761,G6762);
  nand GNAME2443(G2443,G36,G35);
  nand GNAME2444(G2444,G788,G2443);
  nand GNAME2445(G2445,G1200,G36);
  nand GNAME2446(G2446,G2444,G1203);
  nand GNAME2447(G2447,G2445,G2446);
  nand GNAME2448(G2448,G2447,G21392);
  nand GNAME2449(G2449,G2442,G21390);
  nand GNAME2450(G2450,G6744,G6745);
  or GNAME2451(G2451,G788,G33);
  nand GNAME2452(G2452,G1195,G35);
  nand GNAME2453(G2453,G788,G21390);
  nand GNAME2454(G2454,G2453,G2441);
  nand GNAME2455(G2455,G1194,G2451);
  nand GNAME2456(G2456,G2455,G21390);
  or GNAME2457(G2457,G1589,G34);
  nor GNAME2458(G2458,G21391,G1197);
  or GNAME2459(G2459,G2458,G1201);
  not GNAME2460(G2460,G1246);
  nand GNAME2461(G2461,G1216,G21431);
  nand GNAME2462(G2462,G1218,G21439);
  nand GNAME2463(G2463,G1220,G21447);
  nand GNAME2464(G2464,G1222,G21455);
  nand GNAME2465(G2465,G1224,G21463);
  nand GNAME2466(G2466,G1225,G21471);
  nand GNAME2467(G2467,G1226,G21479);
  nand GNAME2468(G2468,G1227,G21487);
  nand GNAME2469(G2469,G1229,G21495);
  nand GNAME2470(G2470,G1230,G21503);
  nand GNAME2471(G2471,G1231,G21511);
  nand GNAME2472(G2472,G1232,G21519);
  nand GNAME2473(G2473,G1234,G21527);
  nand GNAME2474(G2474,G1235,G21535);
  nand GNAME2475(G2475,G1236,G21543);
  nand GNAME2476(G2476,G1237,G21551);
  not GNAME2477(G2477,G1242);
  nand GNAME2478(G2478,G1216,G21432);
  nand GNAME2479(G2479,G1218,G21440);
  nand GNAME2480(G2480,G1220,G21448);
  nand GNAME2481(G2481,G1222,G21456);
  nand GNAME2482(G2482,G1224,G21464);
  nand GNAME2483(G2483,G1225,G21472);
  nand GNAME2484(G2484,G1226,G21480);
  nand GNAME2485(G2485,G1227,G21488);
  nand GNAME2486(G2486,G1229,G21496);
  nand GNAME2487(G2487,G1230,G21504);
  nand GNAME2488(G2488,G1231,G21512);
  nand GNAME2489(G2489,G1232,G21520);
  nand GNAME2490(G2490,G1234,G21528);
  nand GNAME2491(G2491,G1235,G21536);
  nand GNAME2492(G2492,G1236,G21544);
  nand GNAME2493(G2493,G1237,G21552);
  not GNAME2494(G2494,G1192);
  nand GNAME2495(G2495,G1216,G21436);
  nand GNAME2496(G2496,G1218,G21444);
  nand GNAME2497(G2497,G1220,G21452);
  nand GNAME2498(G2498,G1222,G21460);
  nand GNAME2499(G2499,G1224,G21468);
  nand GNAME2500(G2500,G1225,G21476);
  nand GNAME2501(G2501,G1226,G21484);
  nand GNAME2502(G2502,G1227,G21492);
  nand GNAME2503(G2503,G1229,G21500);
  nand GNAME2504(G2504,G1230,G21508);
  nand GNAME2505(G2505,G1231,G21516);
  nand GNAME2506(G2506,G1232,G21524);
  nand GNAME2507(G2507,G1234,G21532);
  nand GNAME2508(G2508,G1235,G21540);
  nand GNAME2509(G2509,G1236,G21548);
  nand GNAME2510(G2510,G1237,G21556);
  not GNAME2511(G2511,G1248);
  nand GNAME2512(G2512,G1216,G21430);
  nand GNAME2513(G2513,G1218,G21438);
  nand GNAME2514(G2514,G1220,G21446);
  nand GNAME2515(G2515,G1222,G21454);
  nand GNAME2516(G2516,G1224,G21462);
  nand GNAME2517(G2517,G1225,G21470);
  nand GNAME2518(G2518,G1226,G21478);
  nand GNAME2519(G2519,G1227,G21486);
  nand GNAME2520(G2520,G1229,G21494);
  nand GNAME2521(G2521,G1230,G21502);
  nand GNAME2522(G2522,G1231,G21510);
  nand GNAME2523(G2523,G1232,G21518);
  nand GNAME2524(G2524,G1234,G21526);
  nand GNAME2525(G2525,G1235,G21534);
  nand GNAME2526(G2526,G1236,G21542);
  nand GNAME2527(G2527,G1237,G21550);
  not GNAME2528(G2528,G1239);
  nand GNAME2529(G2529,G1216,G21435);
  nand GNAME2530(G2530,G1218,G21443);
  nand GNAME2531(G2531,G1220,G21451);
  nand GNAME2532(G2532,G1222,G21459);
  nand GNAME2533(G2533,G1224,G21467);
  nand GNAME2534(G2534,G1225,G21475);
  nand GNAME2535(G2535,G1226,G21483);
  nand GNAME2536(G2536,G1227,G21491);
  nand GNAME2537(G2537,G1229,G21499);
  nand GNAME2538(G2538,G1230,G21507);
  nand GNAME2539(G2539,G1231,G21515);
  nand GNAME2540(G2540,G1232,G21523);
  nand GNAME2541(G2541,G1234,G21531);
  nand GNAME2542(G2542,G1235,G21539);
  nand GNAME2543(G2543,G1236,G21547);
  nand GNAME2544(G2544,G1237,G21555);
  not GNAME2545(G2545,G1238);
  nand GNAME2546(G2546,G1216,G21433);
  nand GNAME2547(G2547,G1218,G21441);
  nand GNAME2548(G2548,G1220,G21449);
  nand GNAME2549(G2549,G1222,G21457);
  nand GNAME2550(G2550,G1224,G21465);
  nand GNAME2551(G2551,G1225,G21473);
  nand GNAME2552(G2552,G1226,G21481);
  nand GNAME2553(G2553,G1227,G21489);
  nand GNAME2554(G2554,G1229,G21497);
  nand GNAME2555(G2555,G1230,G21505);
  nand GNAME2556(G2556,G1231,G21513);
  nand GNAME2557(G2557,G1232,G21521);
  nand GNAME2558(G2558,G1234,G21529);
  nand GNAME2559(G2559,G1235,G21537);
  nand GNAME2560(G2560,G1236,G21545);
  nand GNAME2561(G2561,G1237,G21553);
  not GNAME2562(G2562,G1249);
  nand GNAME2563(G2563,G1216,G21429);
  nand GNAME2564(G2564,G1218,G21437);
  nand GNAME2565(G2565,G1220,G21445);
  nand GNAME2566(G2566,G1222,G21453);
  nand GNAME2567(G2567,G1224,G21461);
  nand GNAME2568(G2568,G1225,G21469);
  nand GNAME2569(G2569,G1226,G21477);
  nand GNAME2570(G2570,G1227,G21485);
  nand GNAME2571(G2571,G1229,G21493);
  nand GNAME2572(G2572,G1230,G21501);
  nand GNAME2573(G2573,G1231,G21509);
  nand GNAME2574(G2574,G1232,G21517);
  nand GNAME2575(G2575,G1234,G21525);
  nand GNAME2576(G2576,G1235,G21533);
  nand GNAME2577(G2577,G1236,G21541);
  nand GNAME2578(G2578,G1237,G21549);
  not GNAME2579(G2579,G1252);
  nand GNAME2580(G2580,G1216,G21434);
  nand GNAME2581(G2581,G1218,G21442);
  nand GNAME2582(G2582,G1220,G21450);
  nand GNAME2583(G2583,G1222,G21458);
  nand GNAME2584(G2584,G1224,G21466);
  nand GNAME2585(G2585,G1225,G21474);
  nand GNAME2586(G2586,G1226,G21482);
  nand GNAME2587(G2587,G1227,G21490);
  nand GNAME2588(G2588,G1229,G21498);
  nand GNAME2589(G2589,G1230,G21506);
  nand GNAME2590(G2590,G1231,G21514);
  nand GNAME2591(G2591,G1232,G21522);
  nand GNAME2592(G2592,G1234,G21530);
  nand GNAME2593(G2593,G1235,G21538);
  nand GNAME2594(G2594,G1236,G21546);
  nand GNAME2595(G2595,G1237,G21554);
  not GNAME2596(G2596,G1240);
  or GNAME2597(G2597,G21428,G21427);
  not GNAME2598(G2598,G1501);
  nand GNAME2599(G2599,G2511,G1251);
  not GNAME2600(G2600,G1253);
  nand GNAME2601(G2601,G1502,G1238);
  nand GNAME2602(G2602,G1253,G2601,G2477);
  nand GNAME2603(G2603,G1238,G2596);
  nand GNAME2604(G2604,G1282,G2603);
  nand GNAME2605(G2605,G2602,G2596);
  nand GNAME2606(G2606,G2596,G1202,G1238);
  nand GNAME2607(G2607,G1204,G1255);
  not GNAME2608(G2608,G682);
  not GNAME2609(G2609,G1263);
  or GNAME2610(G2610,G1263,G2320,G1503);
  nor GNAME2611(G2611,G21795,G21796);
  not GNAME2612(G2612,G1268);
  nand GNAME2613(G2613,G1272,G2612);
  or GNAME2614(G2614,G1247,G1245,G1246);
  not GNAME2615(G2615,G1273);
  nand GNAME2616(G2616,G1275,G1202,G21427);
  nand GNAME2617(G2617,G1269,G1277);
  nand GNAME2618(G2618,G1202,G1280);
  nand GNAME2619(G2619,G2618,G2332);
  nand GNAME2620(G2620,G2341,G1271);
  nand GNAME2621(G2621,G21428,G1271,G2619);
  nand GNAME2622(G2622,G2620,G21427);
  nand GNAME2623(G2623,G7326,G21425,G1281);
  nand GNAME2624(G2624,G1273,G7326);
  nand GNAME2625(G2625,G1269,G2623);
  nand GNAME2626(G2626,G1268,G1283);
  nand GNAME2627(G2627,G2626,G2624,G2625);
  nand GNAME2628(G2628,G2278,G21563);
  not GNAME2629(G2629,G1433);
  nand GNAME2630(G2630,G1299,G21558);
  nand GNAME2631(G2631,G21563,G1292);
  nand GNAME2632(G2632,G1209,G1433);
  nand GNAME2633(G2633,G1273,G6788,G6789);
  not GNAME2634(G2634,G1304);
  nand GNAME2635(G2635,G21565,G21566);
  and GNAME2636(G2636,G2635,G21564);
  not GNAME2637(G2637,G1388);
  nand GNAME2638(G2638,G1299,G21559);
  nand GNAME2639(G2639,G21564,G1292);
  nand GNAME2640(G2640,G1209,G1388);
  not GNAME2641(G2641,G1309);
  not GNAME2642(G2642,G1363);
  nand GNAME2643(G2643,G1299,G21560);
  nand GNAME2644(G2644,G21565,G1292);
  nand GNAME2645(G2645,G1209,G1363);
  not GNAME2646(G2646,G1305);
  nor GNAME2647(G2647,G21427,G1264);
  not GNAME2648(G2648,G1302);
  nand GNAME2649(G2649,G1299,G21561);
  not GNAME2650(G2650,G1301);
  not GNAME2651(G2651,G1306);
  nand GNAME2652(G2652,G1305,G1306);
  nand GNAME2653(G2653,G2652,G2634);
  nand GNAME2654(G2654,G2651,G2646);
  and GNAME2655(G2655,G1296,G2459,G1238);
  not GNAME2656(G2656,G1298);
  not GNAME2657(G2657,G1312);
  or GNAME2658(G2658,G1209,G1297);
  nand GNAME2659(G2659,G2656,G2657,G2658);
  nand GNAME2660(G2660,G2659,G21558);
  nand GNAME2661(G2661,G1209,G6804);
  nand GNAME2662(G2662,G1304,G2654);
  nand GNAME2663(G2663,G2641,G2662,G2652);
  nand GNAME2664(G2664,G2659,G21559);
  nand GNAME2665(G2665,G1209,G2259);
  not GNAME2666(G2666,G1314);
  nand GNAME2667(G2667,G2659,G21560);
  nand GNAME2668(G2668,G1209,G1727);
  not GNAME2669(G2669,G1307);
  nand GNAME2670(G2670,G2650,G2648);
  nand GNAME2671(G2671,G2659,G21561);
  nand GNAME2672(G2672,G1209,G2258);
  not GNAME2673(G2673,G1308);
  nand GNAME2674(G2674,G1298,G2673);
  nand GNAME2675(G2675,G2674,G2669);
  nand GNAME2676(G2676,G1308,G2656);
  not GNAME2677(G2677,G1311);
  nand GNAME2678(G2678,G2657,G1311);
  nand GNAME2679(G2679,G1314,G2678);
  nand GNAME2680(G2680,G2677,G1312);
  nand GNAME2681(G2681,G1312,G2666);
  nand GNAME2682(G2682,G2657,G1314);
  nand GNAME2683(G2683,G2681,G2682);
  nand GNAME2684(G2684,G1296,G1313);
  nand GNAME2685(G2685,G6810,G1320);
  nand GNAME2686(G2686,G25,G1322);
  nand GNAME2687(G2687,G9,G2286);
  nand GNAME2688(G2688,G2687,G2685,G2686);
  nand GNAME2689(G2689,G7326,G1291);
  not GNAME2690(G2690,G1531);
  nand GNAME2691(G2691,G1323,G21426);
  nand GNAME2692(G2692,G2691,G2317);
  nand GNAME2693(G2693,G2294,G2692);
  nand GNAME2694(G2694,G2693,G1531);
  or GNAME2695(G2695,G2298,G1321);
  nand GNAME2696(G2696,G21426,G2286);
  nand GNAME2697(G2697,G2695,G2696);
  nand GNAME2698(G2698,G1252,G1281);
  nand GNAME2699(G2699,G21426,G25);
  nand GNAME2700(G2700,G2698,G2699);
  nand GNAME2701(G2701,G6810,G1295);
  nand GNAME2702(G2702,G2688,G1324);
  nand GNAME2703(G2703,G1325,G1326);
  nand GNAME2704(G2704,G1294,G1327);
  nand GNAME2705(G2705,G2697,G1328);
  nand GNAME2706(G2706,G2694,G21429);
  nand GNAME2707(G2707,G6813,G1320);
  nand GNAME2708(G2708,G1322,G26);
  nand GNAME2709(G2709,G2286,G10);
  nand GNAME2710(G2710,G2709,G2707,G2708);
  nand GNAME2711(G2711,G1239,G1281);
  nand GNAME2712(G2712,G21426,G26);
  nand GNAME2713(G2713,G2711,G2712);
  nand GNAME2714(G2714,G6813,G1295);
  nand GNAME2715(G2715,G2710,G1324);
  nand GNAME2716(G2716,G1326,G1329);
  nand GNAME2717(G2717,G1294,G1330);
  nand GNAME2718(G2718,G2697,G1331);
  nand GNAME2719(G2719,G2694,G21430);
  nand GNAME2720(G2720,G6816,G1320);
  nand GNAME2721(G2721,G1322,G27);
  nand GNAME2722(G2722,G2286,G11);
  nand GNAME2723(G2723,G2722,G2720,G2721);
  nand GNAME2724(G2724,G1242,G1281);
  nand GNAME2725(G2725,G21426,G27);
  nand GNAME2726(G2726,G2724,G2725);
  nand GNAME2727(G2727,G6816,G1295);
  nand GNAME2728(G2728,G2723,G1324);
  nand GNAME2729(G2729,G1326,G1332);
  nand GNAME2730(G2730,G1294,G1333);
  nand GNAME2731(G2731,G2697,G1334);
  nand GNAME2732(G2732,G2694,G21431);
  nand GNAME2733(G2733,G6819,G1320);
  nand GNAME2734(G2734,G1322,G28);
  nand GNAME2735(G2735,G2286,G12);
  nand GNAME2736(G2736,G2735,G2733,G2734);
  nand GNAME2737(G2737,G1192,G1281);
  nand GNAME2738(G2738,G21426,G28);
  nand GNAME2739(G2739,G2737,G2738);
  nand GNAME2740(G2740,G6819,G1295);
  nand GNAME2741(G2741,G2736,G1324);
  nand GNAME2742(G2742,G1326,G1335);
  nand GNAME2743(G2743,G1294,G1336);
  nand GNAME2744(G2744,G2697,G1337);
  nand GNAME2745(G2745,G2694,G21432);
  nand GNAME2746(G2746,G6822,G1320);
  nand GNAME2747(G2747,G1322,G29);
  nand GNAME2748(G2748,G2286,G13);
  nand GNAME2749(G2749,G2748,G2746,G2747);
  nand GNAME2750(G2750,G1249,G1281);
  nand GNAME2751(G2751,G21426,G29);
  nand GNAME2752(G2752,G2750,G2751);
  nand GNAME2753(G2753,G6822,G1295);
  nand GNAME2754(G2754,G2749,G1324);
  nand GNAME2755(G2755,G1326,G1338);
  nand GNAME2756(G2756,G1294,G1339);
  nand GNAME2757(G2757,G2697,G1340);
  nand GNAME2758(G2758,G2694,G21433);
  nand GNAME2759(G2759,G6825,G1320);
  nand GNAME2760(G2760,G1322,G30);
  nand GNAME2761(G2761,G2286,G14);
  nand GNAME2762(G2762,G2761,G2759,G2760);
  nand GNAME2763(G2763,G1240,G1281);
  nand GNAME2764(G2764,G21426,G30);
  nand GNAME2765(G2765,G2763,G2764);
  nand GNAME2766(G2766,G6825,G1295);
  nand GNAME2767(G2767,G2762,G1324);
  nand GNAME2768(G2768,G1326,G1341);
  nand GNAME2769(G2769,G1294,G1342);
  nand GNAME2770(G2770,G2697,G1343);
  nand GNAME2771(G2771,G2694,G21434);
  nand GNAME2772(G2772,G6828,G1320);
  nand GNAME2773(G2773,G1322,G31);
  nand GNAME2774(G2774,G2286,G15);
  nand GNAME2775(G2775,G2774,G2772,G2773);
  nand GNAME2776(G2776,G1238,G1281);
  nand GNAME2777(G2777,G21426,G31);
  nand GNAME2778(G2778,G2776,G2777);
  nand GNAME2779(G2779,G6828,G1295);
  nand GNAME2780(G2780,G2775,G1324);
  nand GNAME2781(G2781,G1326,G1344);
  nand GNAME2782(G2782,G1294,G1345);
  nand GNAME2783(G2783,G2697,G1346);
  nand GNAME2784(G2784,G2694,G21435);
  nand GNAME2785(G2785,G6831,G1320);
  nand GNAME2786(G2786,G1322,G32);
  nand GNAME2787(G2787,G2286,G16);
  nand GNAME2788(G2788,G2787,G2785,G2786);
  nand GNAME2789(G2789,G1248,G1281);
  nand GNAME2790(G2790,G21426,G32);
  nand GNAME2791(G2791,G2789,G2790);
  nand GNAME2792(G2792,G6831,G1295);
  nand GNAME2793(G2793,G2788,G1324);
  nand GNAME2794(G2794,G1326,G1347);
  nand GNAME2795(G2795,G1294,G1348);
  nand GNAME2796(G2796,G2697,G1349);
  nand GNAME2797(G2797,G2694,G21436);
  nand GNAME2798(G2798,G6834,G1357);
  nand GNAME2799(G2799,G25,G1359);
  nand GNAME2800(G2800,G9,G2285);
  nand GNAME2801(G2801,G2800,G2798,G2799);
  nand GNAME2802(G2802,G1360,G21426);
  nand GNAME2803(G2803,G2802,G2317);
  nand GNAME2804(G2804,G1353,G2803);
  nand GNAME2805(G2805,G2804,G1531);
  or GNAME2806(G2806,G2298,G1358);
  nand GNAME2807(G2807,G21426,G2285);
  nand GNAME2808(G2808,G2806,G2807);
  nand GNAME2809(G2809,G6834,G1354);
  nand GNAME2810(G2810,G2801,G1361);
  nand GNAME2811(G2811,G1325,G1362);
  nand GNAME2812(G2812,G1327,G2293);
  nand GNAME2813(G2813,G2808,G1328);
  nand GNAME2814(G2814,G2805,G21437);
  nand GNAME2815(G2815,G6837,G1357);
  nand GNAME2816(G2816,G26,G1359);
  nand GNAME2817(G2817,G10,G2285);
  nand GNAME2818(G2818,G2817,G2815,G2816);
  nand GNAME2819(G2819,G6837,G1354);
  nand GNAME2820(G2820,G2818,G1361);
  nand GNAME2821(G2821,G1329,G1362);
  nand GNAME2822(G2822,G1330,G2293);
  nand GNAME2823(G2823,G2808,G1331);
  nand GNAME2824(G2824,G2805,G21438);
  nand GNAME2825(G2825,G6840,G1357);
  nand GNAME2826(G2826,G27,G1359);
  nand GNAME2827(G2827,G11,G2285);
  nand GNAME2828(G2828,G2827,G2825,G2826);
  nand GNAME2829(G2829,G6840,G1354);
  nand GNAME2830(G2830,G2828,G1361);
  nand GNAME2831(G2831,G1332,G1362);
  nand GNAME2832(G2832,G1333,G2293);
  nand GNAME2833(G2833,G2808,G1334);
  nand GNAME2834(G2834,G2805,G21439);
  nand GNAME2835(G2835,G6843,G1357);
  nand GNAME2836(G2836,G28,G1359);
  nand GNAME2837(G2837,G12,G2285);
  nand GNAME2838(G2838,G2837,G2835,G2836);
  nand GNAME2839(G2839,G6843,G1354);
  nand GNAME2840(G2840,G2838,G1361);
  nand GNAME2841(G2841,G1335,G1362);
  nand GNAME2842(G2842,G1336,G2293);
  nand GNAME2843(G2843,G2808,G1337);
  nand GNAME2844(G2844,G2805,G21440);
  nand GNAME2845(G2845,G6846,G1357);
  nand GNAME2846(G2846,G29,G1359);
  nand GNAME2847(G2847,G13,G2285);
  nand GNAME2848(G2848,G2847,G2845,G2846);
  nand GNAME2849(G2849,G6846,G1354);
  nand GNAME2850(G2850,G2848,G1361);
  nand GNAME2851(G2851,G1338,G1362);
  nand GNAME2852(G2852,G1339,G2293);
  nand GNAME2853(G2853,G2808,G1340);
  nand GNAME2854(G2854,G2805,G21441);
  nand GNAME2855(G2855,G6849,G1357);
  nand GNAME2856(G2856,G30,G1359);
  nand GNAME2857(G2857,G14,G2285);
  nand GNAME2858(G2858,G2857,G2855,G2856);
  nand GNAME2859(G2859,G6849,G1354);
  nand GNAME2860(G2860,G2858,G1361);
  nand GNAME2861(G2861,G1341,G1362);
  nand GNAME2862(G2862,G1342,G2293);
  nand GNAME2863(G2863,G2808,G1343);
  nand GNAME2864(G2864,G2805,G21442);
  nand GNAME2865(G2865,G6852,G1357);
  nand GNAME2866(G2866,G31,G1359);
  nand GNAME2867(G2867,G15,G2285);
  nand GNAME2868(G2868,G2867,G2865,G2866);
  nand GNAME2869(G2869,G6852,G1354);
  nand GNAME2870(G2870,G2868,G1361);
  nand GNAME2871(G2871,G1344,G1362);
  nand GNAME2872(G2872,G1345,G2293);
  nand GNAME2873(G2873,G2808,G1346);
  nand GNAME2874(G2874,G2805,G21443);
  nand GNAME2875(G2875,G6855,G1357);
  nand GNAME2876(G2876,G32,G1359);
  nand GNAME2877(G2877,G16,G2285);
  nand GNAME2878(G2878,G2877,G2875,G2876);
  nand GNAME2879(G2879,G6855,G1354);
  nand GNAME2880(G2880,G2878,G1361);
  nand GNAME2881(G2881,G1347,G1362);
  nand GNAME2882(G2882,G1348,G2293);
  nand GNAME2883(G2883,G2808,G1349);
  nand GNAME2884(G2884,G2805,G21444);
  nand GNAME2885(G2885,G6858,G1371);
  nand GNAME2886(G2886,G25,G1373);
  nand GNAME2887(G2887,G9,G2284);
  nand GNAME2888(G2888,G2887,G2885,G2886);
  nand GNAME2889(G2889,G1374,G21426);
  nand GNAME2890(G2890,G2889,G2317);
  nand GNAME2891(G2891,G1367,G2890);
  nand GNAME2892(G2892,G2891,G1531);
  or GNAME2893(G2893,G2298,G1372);
  nand GNAME2894(G2894,G21426,G2284);
  nand GNAME2895(G2895,G2893,G2894);
  nand GNAME2896(G2896,G6858,G1368);
  nand GNAME2897(G2897,G2888,G1375);
  nand GNAME2898(G2898,G1325,G1376);
  nand GNAME2899(G2899,G1327,G2292);
  nand GNAME2900(G2900,G2895,G1328);
  nand GNAME2901(G2901,G2892,G21445);
  nand GNAME2902(G2902,G6861,G1371);
  nand GNAME2903(G2903,G26,G1373);
  nand GNAME2904(G2904,G10,G2284);
  nand GNAME2905(G2905,G2904,G2902,G2903);
  nand GNAME2906(G2906,G6861,G1368);
  nand GNAME2907(G2907,G2905,G1375);
  nand GNAME2908(G2908,G1329,G1376);
  nand GNAME2909(G2909,G1330,G2292);
  nand GNAME2910(G2910,G2895,G1331);
  nand GNAME2911(G2911,G2892,G21446);
  nand GNAME2912(G2912,G6864,G1371);
  nand GNAME2913(G2913,G27,G1373);
  nand GNAME2914(G2914,G11,G2284);
  nand GNAME2915(G2915,G2914,G2912,G2913);
  nand GNAME2916(G2916,G6864,G1368);
  nand GNAME2917(G2917,G2915,G1375);
  nand GNAME2918(G2918,G1332,G1376);
  nand GNAME2919(G2919,G1333,G2292);
  nand GNAME2920(G2920,G2895,G1334);
  nand GNAME2921(G2921,G2892,G21447);
  nand GNAME2922(G2922,G6867,G1371);
  nand GNAME2923(G2923,G28,G1373);
  nand GNAME2924(G2924,G12,G2284);
  nand GNAME2925(G2925,G2924,G2922,G2923);
  nand GNAME2926(G2926,G6867,G1368);
  nand GNAME2927(G2927,G2925,G1375);
  nand GNAME2928(G2928,G1335,G1376);
  nand GNAME2929(G2929,G1336,G2292);
  nand GNAME2930(G2930,G2895,G1337);
  nand GNAME2931(G2931,G2892,G21448);
  nand GNAME2932(G2932,G6870,G1371);
  nand GNAME2933(G2933,G29,G1373);
  nand GNAME2934(G2934,G13,G2284);
  nand GNAME2935(G2935,G2934,G2932,G2933);
  nand GNAME2936(G2936,G6870,G1368);
  nand GNAME2937(G2937,G2935,G1375);
  nand GNAME2938(G2938,G1338,G1376);
  nand GNAME2939(G2939,G1339,G2292);
  nand GNAME2940(G2940,G2895,G1340);
  nand GNAME2941(G2941,G2892,G21449);
  nand GNAME2942(G2942,G6873,G1371);
  nand GNAME2943(G2943,G30,G1373);
  nand GNAME2944(G2944,G14,G2284);
  nand GNAME2945(G2945,G2944,G2942,G2943);
  nand GNAME2946(G2946,G6873,G1368);
  nand GNAME2947(G2947,G2945,G1375);
  nand GNAME2948(G2948,G1341,G1376);
  nand GNAME2949(G2949,G1342,G2292);
  nand GNAME2950(G2950,G2895,G1343);
  nand GNAME2951(G2951,G2892,G21450);
  nand GNAME2952(G2952,G6876,G1371);
  nand GNAME2953(G2953,G31,G1373);
  nand GNAME2954(G2954,G15,G2284);
  nand GNAME2955(G2955,G2954,G2952,G2953);
  nand GNAME2956(G2956,G6876,G1368);
  nand GNAME2957(G2957,G2955,G1375);
  nand GNAME2958(G2958,G1344,G1376);
  nand GNAME2959(G2959,G1345,G2292);
  nand GNAME2960(G2960,G2895,G1346);
  nand GNAME2961(G2961,G2892,G21451);
  nand GNAME2962(G2962,G6879,G1371);
  nand GNAME2963(G2963,G32,G1373);
  nand GNAME2964(G2964,G16,G2284);
  nand GNAME2965(G2965,G2964,G2962,G2963);
  nand GNAME2966(G2966,G6879,G1368);
  nand GNAME2967(G2967,G2965,G1375);
  nand GNAME2968(G2968,G1347,G1376);
  nand GNAME2969(G2969,G1348,G2292);
  nand GNAME2970(G2970,G2895,G1349);
  nand GNAME2971(G2971,G2892,G21452);
  nand GNAME2972(G2972,G6882,G1382);
  nand GNAME2973(G2973,G25,G1384);
  nand GNAME2974(G2974,G9,G2283);
  nand GNAME2975(G2975,G2974,G2972,G2973);
  nand GNAME2976(G2976,G1385,G21426);
  nand GNAME2977(G2977,G2976,G2317);
  nand GNAME2978(G2978,G1379,G2977);
  nand GNAME2979(G2979,G2978,G1531);
  or GNAME2980(G2980,G2298,G1383);
  nand GNAME2981(G2981,G21426,G2283);
  nand GNAME2982(G2982,G2980,G2981);
  nand GNAME2983(G2983,G6882,G1380);
  nand GNAME2984(G2984,G2975,G1386);
  nand GNAME2985(G2985,G1325,G1387);
  nand GNAME2986(G2986,G1327,G2291);
  nand GNAME2987(G2987,G2982,G1328);
  nand GNAME2988(G2988,G2979,G21453);
  nand GNAME2989(G2989,G6885,G1382);
  nand GNAME2990(G2990,G26,G1384);
  nand GNAME2991(G2991,G10,G2283);
  nand GNAME2992(G2992,G2991,G2989,G2990);
  nand GNAME2993(G2993,G6885,G1380);
  nand GNAME2994(G2994,G2992,G1386);
  nand GNAME2995(G2995,G1329,G1387);
  nand GNAME2996(G2996,G1330,G2291);
  nand GNAME2997(G2997,G2982,G1331);
  nand GNAME2998(G2998,G2979,G21454);
  nand GNAME2999(G2999,G6888,G1382);
  nand GNAME3000(G3000,G27,G1384);
  nand GNAME3001(G3001,G11,G2283);
  nand GNAME3002(G3002,G3001,G2999,G3000);
  nand GNAME3003(G3003,G6888,G1380);
  nand GNAME3004(G3004,G3002,G1386);
  nand GNAME3005(G3005,G1332,G1387);
  nand GNAME3006(G3006,G1333,G2291);
  nand GNAME3007(G3007,G2982,G1334);
  nand GNAME3008(G3008,G2979,G21455);
  nand GNAME3009(G3009,G6891,G1382);
  nand GNAME3010(G3010,G28,G1384);
  nand GNAME3011(G3011,G12,G2283);
  nand GNAME3012(G3012,G3011,G3009,G3010);
  nand GNAME3013(G3013,G6891,G1380);
  nand GNAME3014(G3014,G3012,G1386);
  nand GNAME3015(G3015,G1335,G1387);
  nand GNAME3016(G3016,G1336,G2291);
  nand GNAME3017(G3017,G2982,G1337);
  nand GNAME3018(G3018,G2979,G21456);
  nand GNAME3019(G3019,G6894,G1382);
  nand GNAME3020(G3020,G29,G1384);
  nand GNAME3021(G3021,G13,G2283);
  nand GNAME3022(G3022,G3021,G3019,G3020);
  nand GNAME3023(G3023,G6894,G1380);
  nand GNAME3024(G3024,G3022,G1386);
  nand GNAME3025(G3025,G1338,G1387);
  nand GNAME3026(G3026,G1339,G2291);
  nand GNAME3027(G3027,G2982,G1340);
  nand GNAME3028(G3028,G2979,G21457);
  nand GNAME3029(G3029,G6897,G1382);
  nand GNAME3030(G3030,G30,G1384);
  nand GNAME3031(G3031,G14,G2283);
  nand GNAME3032(G3032,G3031,G3029,G3030);
  nand GNAME3033(G3033,G6897,G1380);
  nand GNAME3034(G3034,G3032,G1386);
  nand GNAME3035(G3035,G1341,G1387);
  nand GNAME3036(G3036,G1342,G2291);
  nand GNAME3037(G3037,G2982,G1343);
  nand GNAME3038(G3038,G2979,G21458);
  nand GNAME3039(G3039,G6900,G1382);
  nand GNAME3040(G3040,G31,G1384);
  nand GNAME3041(G3041,G15,G2283);
  nand GNAME3042(G3042,G3041,G3039,G3040);
  nand GNAME3043(G3043,G6900,G1380);
  nand GNAME3044(G3044,G3042,G1386);
  nand GNAME3045(G3045,G1344,G1387);
  nand GNAME3046(G3046,G1345,G2291);
  nand GNAME3047(G3047,G2982,G1346);
  nand GNAME3048(G3048,G2979,G21459);
  nand GNAME3049(G3049,G6903,G1382);
  nand GNAME3050(G3050,G32,G1384);
  nand GNAME3051(G3051,G16,G2283);
  nand GNAME3052(G3052,G3051,G3049,G3050);
  nand GNAME3053(G3053,G6903,G1380);
  nand GNAME3054(G3054,G3052,G1386);
  nand GNAME3055(G3055,G1347,G1387);
  nand GNAME3056(G3056,G1348,G2291);
  nand GNAME3057(G3057,G2982,G1349);
  nand GNAME3058(G3058,G2979,G21460);
  nand GNAME3059(G3059,G6906,G1395);
  nand GNAME3060(G3060,G25,G1397);
  nand GNAME3061(G3061,G9,G2282);
  nand GNAME3062(G3062,G3061,G3059,G3060);
  nand GNAME3063(G3063,G1398,G21426);
  nand GNAME3064(G3064,G3063,G2317);
  nand GNAME3065(G3065,G1391,G3064);
  nand GNAME3066(G3066,G3065,G1531);
  or GNAME3067(G3067,G2298,G1396);
  nand GNAME3068(G3068,G21426,G2282);
  nand GNAME3069(G3069,G3067,G3068);
  nand GNAME3070(G3070,G6906,G1392);
  nand GNAME3071(G3071,G3062,G1399);
  nand GNAME3072(G3072,G1325,G1400);
  nand GNAME3073(G3073,G1327,G2290);
  nand GNAME3074(G3074,G3069,G1328);
  nand GNAME3075(G3075,G3066,G21461);
  nand GNAME3076(G3076,G6909,G1395);
  nand GNAME3077(G3077,G26,G1397);
  nand GNAME3078(G3078,G10,G2282);
  nand GNAME3079(G3079,G3078,G3076,G3077);
  nand GNAME3080(G3080,G6909,G1392);
  nand GNAME3081(G3081,G3079,G1399);
  nand GNAME3082(G3082,G1329,G1400);
  nand GNAME3083(G3083,G1330,G2290);
  nand GNAME3084(G3084,G3069,G1331);
  nand GNAME3085(G3085,G3066,G21462);
  nand GNAME3086(G3086,G6912,G1395);
  nand GNAME3087(G3087,G27,G1397);
  nand GNAME3088(G3088,G11,G2282);
  nand GNAME3089(G3089,G3088,G3086,G3087);
  nand GNAME3090(G3090,G6912,G1392);
  nand GNAME3091(G3091,G3089,G1399);
  nand GNAME3092(G3092,G1332,G1400);
  nand GNAME3093(G3093,G1333,G2290);
  nand GNAME3094(G3094,G3069,G1334);
  nand GNAME3095(G3095,G3066,G21463);
  nand GNAME3096(G3096,G6915,G1395);
  nand GNAME3097(G3097,G28,G1397);
  nand GNAME3098(G3098,G12,G2282);
  nand GNAME3099(G3099,G3098,G3096,G3097);
  nand GNAME3100(G3100,G6915,G1392);
  nand GNAME3101(G3101,G3099,G1399);
  nand GNAME3102(G3102,G1335,G1400);
  nand GNAME3103(G3103,G1336,G2290);
  nand GNAME3104(G3104,G3069,G1337);
  nand GNAME3105(G3105,G3066,G21464);
  nand GNAME3106(G3106,G6918,G1395);
  nand GNAME3107(G3107,G29,G1397);
  nand GNAME3108(G3108,G13,G2282);
  nand GNAME3109(G3109,G3108,G3106,G3107);
  nand GNAME3110(G3110,G6918,G1392);
  nand GNAME3111(G3111,G3109,G1399);
  nand GNAME3112(G3112,G1338,G1400);
  nand GNAME3113(G3113,G1339,G2290);
  nand GNAME3114(G3114,G3069,G1340);
  nand GNAME3115(G3115,G3066,G21465);
  nand GNAME3116(G3116,G6921,G1395);
  nand GNAME3117(G3117,G30,G1397);
  nand GNAME3118(G3118,G14,G2282);
  nand GNAME3119(G3119,G3118,G3116,G3117);
  nand GNAME3120(G3120,G6921,G1392);
  nand GNAME3121(G3121,G3119,G1399);
  nand GNAME3122(G3122,G1341,G1400);
  nand GNAME3123(G3123,G1342,G2290);
  nand GNAME3124(G3124,G3069,G1343);
  nand GNAME3125(G3125,G3066,G21466);
  nand GNAME3126(G3126,G6924,G1395);
  nand GNAME3127(G3127,G31,G1397);
  nand GNAME3128(G3128,G15,G2282);
  nand GNAME3129(G3129,G3128,G3126,G3127);
  nand GNAME3130(G3130,G6924,G1392);
  nand GNAME3131(G3131,G3129,G1399);
  nand GNAME3132(G3132,G1344,G1400);
  nand GNAME3133(G3133,G1345,G2290);
  nand GNAME3134(G3134,G3069,G1346);
  nand GNAME3135(G3135,G3066,G21467);
  nand GNAME3136(G3136,G6927,G1395);
  nand GNAME3137(G3137,G32,G1397);
  nand GNAME3138(G3138,G16,G2282);
  nand GNAME3139(G3139,G3138,G3136,G3137);
  nand GNAME3140(G3140,G6927,G1392);
  nand GNAME3141(G3141,G3139,G1399);
  nand GNAME3142(G3142,G1347,G1400);
  nand GNAME3143(G3143,G1348,G2290);
  nand GNAME3144(G3144,G3069,G1349);
  nand GNAME3145(G3145,G3066,G21468);
  nand GNAME3146(G3146,G6930,G1406);
  nand GNAME3147(G3147,G25,G1408);
  nand GNAME3148(G3148,G9,G2281);
  nand GNAME3149(G3149,G3148,G3146,G3147);
  nand GNAME3150(G3150,G1409,G21426);
  nand GNAME3151(G3151,G3150,G2317);
  nand GNAME3152(G3152,G1402,G3151);
  nand GNAME3153(G3153,G3152,G1531);
  or GNAME3154(G3154,G2298,G1407);
  nand GNAME3155(G3155,G21426,G2281);
  nand GNAME3156(G3156,G3154,G3155);
  nand GNAME3157(G3157,G6930,G1403);
  nand GNAME3158(G3158,G3149,G1410);
  nand GNAME3159(G3159,G1325,G1411);
  nand GNAME3160(G3160,G1327,G2289);
  nand GNAME3161(G3161,G3156,G1328);
  nand GNAME3162(G3162,G3153,G21469);
  nand GNAME3163(G3163,G6933,G1406);
  nand GNAME3164(G3164,G26,G1408);
  nand GNAME3165(G3165,G10,G2281);
  nand GNAME3166(G3166,G3165,G3163,G3164);
  nand GNAME3167(G3167,G6933,G1403);
  nand GNAME3168(G3168,G3166,G1410);
  nand GNAME3169(G3169,G1329,G1411);
  nand GNAME3170(G3170,G1330,G2289);
  nand GNAME3171(G3171,G3156,G1331);
  nand GNAME3172(G3172,G3153,G21470);
  nand GNAME3173(G3173,G6936,G1406);
  nand GNAME3174(G3174,G27,G1408);
  nand GNAME3175(G3175,G11,G2281);
  nand GNAME3176(G3176,G3175,G3173,G3174);
  nand GNAME3177(G3177,G6936,G1403);
  nand GNAME3178(G3178,G3176,G1410);
  nand GNAME3179(G3179,G1332,G1411);
  nand GNAME3180(G3180,G1333,G2289);
  nand GNAME3181(G3181,G3156,G1334);
  nand GNAME3182(G3182,G3153,G21471);
  nand GNAME3183(G3183,G6939,G1406);
  nand GNAME3184(G3184,G28,G1408);
  nand GNAME3185(G3185,G12,G2281);
  nand GNAME3186(G3186,G3185,G3183,G3184);
  nand GNAME3187(G3187,G6939,G1403);
  nand GNAME3188(G3188,G3186,G1410);
  nand GNAME3189(G3189,G1335,G1411);
  nand GNAME3190(G3190,G1336,G2289);
  nand GNAME3191(G3191,G3156,G1337);
  nand GNAME3192(G3192,G3153,G21472);
  nand GNAME3193(G3193,G6942,G1406);
  nand GNAME3194(G3194,G29,G1408);
  nand GNAME3195(G3195,G13,G2281);
  nand GNAME3196(G3196,G3195,G3193,G3194);
  nand GNAME3197(G3197,G6942,G1403);
  nand GNAME3198(G3198,G3196,G1410);
  nand GNAME3199(G3199,G1338,G1411);
  nand GNAME3200(G3200,G1339,G2289);
  nand GNAME3201(G3201,G3156,G1340);
  nand GNAME3202(G3202,G3153,G21473);
  nand GNAME3203(G3203,G6945,G1406);
  nand GNAME3204(G3204,G30,G1408);
  nand GNAME3205(G3205,G14,G2281);
  nand GNAME3206(G3206,G3205,G3203,G3204);
  nand GNAME3207(G3207,G6945,G1403);
  nand GNAME3208(G3208,G3206,G1410);
  nand GNAME3209(G3209,G1341,G1411);
  nand GNAME3210(G3210,G1342,G2289);
  nand GNAME3211(G3211,G3156,G1343);
  nand GNAME3212(G3212,G3153,G21474);
  nand GNAME3213(G3213,G6948,G1406);
  nand GNAME3214(G3214,G31,G1408);
  nand GNAME3215(G3215,G15,G2281);
  nand GNAME3216(G3216,G3215,G3213,G3214);
  nand GNAME3217(G3217,G6948,G1403);
  nand GNAME3218(G3218,G3216,G1410);
  nand GNAME3219(G3219,G1344,G1411);
  nand GNAME3220(G3220,G1345,G2289);
  nand GNAME3221(G3221,G3156,G1346);
  nand GNAME3222(G3222,G3153,G21475);
  nand GNAME3223(G3223,G6951,G1406);
  nand GNAME3224(G3224,G32,G1408);
  nand GNAME3225(G3225,G16,G2281);
  nand GNAME3226(G3226,G3225,G3223,G3224);
  nand GNAME3227(G3227,G6951,G1403);
  nand GNAME3228(G3228,G3226,G1410);
  nand GNAME3229(G3229,G1347,G1411);
  nand GNAME3230(G3230,G1348,G2289);
  nand GNAME3231(G3231,G3156,G1349);
  nand GNAME3232(G3232,G3153,G21476);
  nand GNAME3233(G3233,G6954,G1416);
  nand GNAME3234(G3234,G25,G1418);
  nand GNAME3235(G3235,G9,G2280);
  nand GNAME3236(G3236,G3235,G3233,G3234);
  nand GNAME3237(G3237,G1419,G21426);
  nand GNAME3238(G3238,G3237,G2317);
  nand GNAME3239(G3239,G1413,G3238);
  nand GNAME3240(G3240,G3239,G1531);
  or GNAME3241(G3241,G2298,G1417);
  nand GNAME3242(G3242,G21426,G2280);
  nand GNAME3243(G3243,G3241,G3242);
  nand GNAME3244(G3244,G6954,G1414);
  nand GNAME3245(G3245,G3236,G1420);
  nand GNAME3246(G3246,G1325,G1421);
  nand GNAME3247(G3247,G1327,G2288);
  nand GNAME3248(G3248,G3243,G1328);
  nand GNAME3249(G3249,G3240,G21477);
  nand GNAME3250(G3250,G6957,G1416);
  nand GNAME3251(G3251,G26,G1418);
  nand GNAME3252(G3252,G10,G2280);
  nand GNAME3253(G3253,G3252,G3250,G3251);
  nand GNAME3254(G3254,G6957,G1414);
  nand GNAME3255(G3255,G3253,G1420);
  nand GNAME3256(G3256,G1329,G1421);
  nand GNAME3257(G3257,G1330,G2288);
  nand GNAME3258(G3258,G3243,G1331);
  nand GNAME3259(G3259,G3240,G21478);
  nand GNAME3260(G3260,G6960,G1416);
  nand GNAME3261(G3261,G27,G1418);
  nand GNAME3262(G3262,G11,G2280);
  nand GNAME3263(G3263,G3262,G3260,G3261);
  nand GNAME3264(G3264,G6960,G1414);
  nand GNAME3265(G3265,G3263,G1420);
  nand GNAME3266(G3266,G1332,G1421);
  nand GNAME3267(G3267,G1333,G2288);
  nand GNAME3268(G3268,G3243,G1334);
  nand GNAME3269(G3269,G3240,G21479);
  nand GNAME3270(G3270,G6963,G1416);
  nand GNAME3271(G3271,G28,G1418);
  nand GNAME3272(G3272,G12,G2280);
  nand GNAME3273(G3273,G3272,G3270,G3271);
  nand GNAME3274(G3274,G6963,G1414);
  nand GNAME3275(G3275,G3273,G1420);
  nand GNAME3276(G3276,G1335,G1421);
  nand GNAME3277(G3277,G1336,G2288);
  nand GNAME3278(G3278,G3243,G1337);
  nand GNAME3279(G3279,G3240,G21480);
  nand GNAME3280(G3280,G6966,G1416);
  nand GNAME3281(G3281,G29,G1418);
  nand GNAME3282(G3282,G13,G2280);
  nand GNAME3283(G3283,G3282,G3280,G3281);
  nand GNAME3284(G3284,G6966,G1414);
  nand GNAME3285(G3285,G3283,G1420);
  nand GNAME3286(G3286,G1338,G1421);
  nand GNAME3287(G3287,G1339,G2288);
  nand GNAME3288(G3288,G3243,G1340);
  nand GNAME3289(G3289,G3240,G21481);
  nand GNAME3290(G3290,G6969,G1416);
  nand GNAME3291(G3291,G30,G1418);
  nand GNAME3292(G3292,G14,G2280);
  nand GNAME3293(G3293,G3292,G3290,G3291);
  nand GNAME3294(G3294,G6969,G1414);
  nand GNAME3295(G3295,G3293,G1420);
  nand GNAME3296(G3296,G1341,G1421);
  nand GNAME3297(G3297,G1342,G2288);
  nand GNAME3298(G3298,G3243,G1343);
  nand GNAME3299(G3299,G3240,G21482);
  nand GNAME3300(G3300,G6972,G1416);
  nand GNAME3301(G3301,G31,G1418);
  nand GNAME3302(G3302,G15,G2280);
  nand GNAME3303(G3303,G3302,G3300,G3301);
  nand GNAME3304(G3304,G6972,G1414);
  nand GNAME3305(G3305,G3303,G1420);
  nand GNAME3306(G3306,G1344,G1421);
  nand GNAME3307(G3307,G1345,G2288);
  nand GNAME3308(G3308,G3243,G1346);
  nand GNAME3309(G3309,G3240,G21483);
  nand GNAME3310(G3310,G6975,G1416);
  nand GNAME3311(G3311,G32,G1418);
  nand GNAME3312(G3312,G16,G2280);
  nand GNAME3313(G3313,G3312,G3310,G3311);
  nand GNAME3314(G3314,G6975,G1414);
  nand GNAME3315(G3315,G3313,G1420);
  nand GNAME3316(G3316,G1347,G1421);
  nand GNAME3317(G3317,G1348,G2288);
  nand GNAME3318(G3318,G3243,G1349);
  nand GNAME3319(G3319,G3240,G21484);
  nand GNAME3320(G3320,G6978,G1426);
  nand GNAME3321(G3321,G25,G1428);
  nand GNAME3322(G3322,G9,G2279);
  nand GNAME3323(G3323,G3322,G3320,G3321);
  nand GNAME3324(G3324,G1429,G21426);
  nand GNAME3325(G3325,G3324,G2317);
  nand GNAME3326(G3326,G1423,G3325);
  nand GNAME3327(G3327,G3326,G1531);
  or GNAME3328(G3328,G2298,G1427);
  nand GNAME3329(G3329,G21426,G2279);
  nand GNAME3330(G3330,G3328,G3329);
  nand GNAME3331(G3331,G6978,G1424);
  nand GNAME3332(G3332,G3323,G1430);
  nand GNAME3333(G3333,G1325,G1431);
  nand GNAME3334(G3334,G1327,G2287);
  nand GNAME3335(G3335,G3330,G1328);
  nand GNAME3336(G3336,G3327,G21485);
  nand GNAME3337(G3337,G6981,G1426);
  nand GNAME3338(G3338,G26,G1428);
  nand GNAME3339(G3339,G10,G2279);
  nand GNAME3340(G3340,G3339,G3337,G3338);
  nand GNAME3341(G3341,G6981,G1424);
  nand GNAME3342(G3342,G3340,G1430);
  nand GNAME3343(G3343,G1329,G1431);
  nand GNAME3344(G3344,G1330,G2287);
  nand GNAME3345(G3345,G3330,G1331);
  nand GNAME3346(G3346,G3327,G21486);
  nand GNAME3347(G3347,G6984,G1426);
  nand GNAME3348(G3348,G27,G1428);
  nand GNAME3349(G3349,G11,G2279);
  nand GNAME3350(G3350,G3349,G3347,G3348);
  nand GNAME3351(G3351,G6984,G1424);
  nand GNAME3352(G3352,G3350,G1430);
  nand GNAME3353(G3353,G1332,G1431);
  nand GNAME3354(G3354,G1333,G2287);
  nand GNAME3355(G3355,G3330,G1334);
  nand GNAME3356(G3356,G3327,G21487);
  nand GNAME3357(G3357,G6987,G1426);
  nand GNAME3358(G3358,G28,G1428);
  nand GNAME3359(G3359,G12,G2279);
  nand GNAME3360(G3360,G3359,G3357,G3358);
  nand GNAME3361(G3361,G6987,G1424);
  nand GNAME3362(G3362,G3360,G1430);
  nand GNAME3363(G3363,G1335,G1431);
  nand GNAME3364(G3364,G1336,G2287);
  nand GNAME3365(G3365,G3330,G1337);
  nand GNAME3366(G3366,G3327,G21488);
  nand GNAME3367(G3367,G6990,G1426);
  nand GNAME3368(G3368,G29,G1428);
  nand GNAME3369(G3369,G13,G2279);
  nand GNAME3370(G3370,G3369,G3367,G3368);
  nand GNAME3371(G3371,G6990,G1424);
  nand GNAME3372(G3372,G3370,G1430);
  nand GNAME3373(G3373,G1338,G1431);
  nand GNAME3374(G3374,G1339,G2287);
  nand GNAME3375(G3375,G3330,G1340);
  nand GNAME3376(G3376,G3327,G21489);
  nand GNAME3377(G3377,G6993,G1426);
  nand GNAME3378(G3378,G30,G1428);
  nand GNAME3379(G3379,G14,G2279);
  nand GNAME3380(G3380,G3379,G3377,G3378);
  nand GNAME3381(G3381,G6993,G1424);
  nand GNAME3382(G3382,G3380,G1430);
  nand GNAME3383(G3383,G1341,G1431);
  nand GNAME3384(G3384,G1342,G2287);
  nand GNAME3385(G3385,G3330,G1343);
  nand GNAME3386(G3386,G3327,G21490);
  nand GNAME3387(G3387,G6996,G1426);
  nand GNAME3388(G3388,G31,G1428);
  nand GNAME3389(G3389,G15,G2279);
  nand GNAME3390(G3390,G3389,G3387,G3388);
  nand GNAME3391(G3391,G6996,G1424);
  nand GNAME3392(G3392,G3390,G1430);
  nand GNAME3393(G3393,G1344,G1431);
  nand GNAME3394(G3394,G1345,G2287);
  nand GNAME3395(G3395,G3330,G1346);
  nand GNAME3396(G3396,G3327,G21491);
  nand GNAME3397(G3397,G6999,G1426);
  nand GNAME3398(G3398,G32,G1428);
  nand GNAME3399(G3399,G16,G2279);
  nand GNAME3400(G3400,G3399,G3397,G3398);
  nand GNAME3401(G3401,G6999,G1424);
  nand GNAME3402(G3402,G3400,G1430);
  nand GNAME3403(G3403,G1347,G1431);
  nand GNAME3404(G3404,G1348,G2287);
  nand GNAME3405(G3405,G3330,G1349);
  nand GNAME3406(G3406,G3327,G21492);
  nand GNAME3407(G3407,G7002,G1436);
  nand GNAME3408(G3408,G25,G1438);
  nand GNAME3409(G3409,G9,G2276);
  nand GNAME3410(G3410,G3409,G3407,G3408);
  nand GNAME3411(G3411,G1439,G21426);
  nand GNAME3412(G3412,G3411,G2317);
  nand GNAME3413(G3413,G2268,G3412);
  nand GNAME3414(G3414,G3413,G1531);
  or GNAME3415(G3415,G2298,G1437);
  nand GNAME3416(G3416,G21426,G2276);
  nand GNAME3417(G3417,G3415,G3416);
  nand GNAME3418(G3418,G3410,G1440);
  nand GNAME3419(G3419,G7002,G1441);
  nand GNAME3420(G3420,G1325,G1442);
  nand GNAME3421(G3421,G1327,G1435);
  nand GNAME3422(G3422,G3417,G1328);
  nand GNAME3423(G3423,G3414,G21493);
  nand GNAME3424(G3424,G7005,G1436);
  nand GNAME3425(G3425,G26,G1438);
  nand GNAME3426(G3426,G10,G2276);
  nand GNAME3427(G3427,G3426,G3424,G3425);
  nand GNAME3428(G3428,G3427,G1440);
  nand GNAME3429(G3429,G7005,G1441);
  nand GNAME3430(G3430,G1329,G1442);
  nand GNAME3431(G3431,G1330,G1435);
  nand GNAME3432(G3432,G3417,G1331);
  nand GNAME3433(G3433,G3414,G21494);
  nand GNAME3434(G3434,G7008,G1436);
  nand GNAME3435(G3435,G27,G1438);
  nand GNAME3436(G3436,G11,G2276);
  nand GNAME3437(G3437,G3436,G3434,G3435);
  nand GNAME3438(G3438,G3437,G1440);
  nand GNAME3439(G3439,G7008,G1441);
  nand GNAME3440(G3440,G1332,G1442);
  nand GNAME3441(G3441,G1333,G1435);
  nand GNAME3442(G3442,G3417,G1334);
  nand GNAME3443(G3443,G3414,G21495);
  nand GNAME3444(G3444,G7011,G1436);
  nand GNAME3445(G3445,G28,G1438);
  nand GNAME3446(G3446,G12,G2276);
  nand GNAME3447(G3447,G3446,G3444,G3445);
  nand GNAME3448(G3448,G3447,G1440);
  nand GNAME3449(G3449,G7011,G1441);
  nand GNAME3450(G3450,G1335,G1442);
  nand GNAME3451(G3451,G1336,G1435);
  nand GNAME3452(G3452,G3417,G1337);
  nand GNAME3453(G3453,G3414,G21496);
  nand GNAME3454(G3454,G7014,G1436);
  nand GNAME3455(G3455,G29,G1438);
  nand GNAME3456(G3456,G13,G2276);
  nand GNAME3457(G3457,G3456,G3454,G3455);
  nand GNAME3458(G3458,G3457,G1440);
  nand GNAME3459(G3459,G7014,G1441);
  nand GNAME3460(G3460,G1338,G1442);
  nand GNAME3461(G3461,G1339,G1435);
  nand GNAME3462(G3462,G3417,G1340);
  nand GNAME3463(G3463,G3414,G21497);
  nand GNAME3464(G3464,G7017,G1436);
  nand GNAME3465(G3465,G30,G1438);
  nand GNAME3466(G3466,G14,G2276);
  nand GNAME3467(G3467,G3466,G3464,G3465);
  nand GNAME3468(G3468,G3467,G1440);
  nand GNAME3469(G3469,G7017,G1441);
  nand GNAME3470(G3470,G1341,G1442);
  nand GNAME3471(G3471,G1342,G1435);
  nand GNAME3472(G3472,G3417,G1343);
  nand GNAME3473(G3473,G3414,G21498);
  nand GNAME3474(G3474,G7020,G1436);
  nand GNAME3475(G3475,G31,G1438);
  nand GNAME3476(G3476,G15,G2276);
  nand GNAME3477(G3477,G3476,G3474,G3475);
  nand GNAME3478(G3478,G3477,G1440);
  nand GNAME3479(G3479,G7020,G1441);
  nand GNAME3480(G3480,G1344,G1442);
  nand GNAME3481(G3481,G1345,G1435);
  nand GNAME3482(G3482,G3417,G1346);
  nand GNAME3483(G3483,G3414,G21499);
  nand GNAME3484(G3484,G7023,G1436);
  nand GNAME3485(G3485,G32,G1438);
  nand GNAME3486(G3486,G16,G2276);
  nand GNAME3487(G3487,G3486,G3484,G3485);
  nand GNAME3488(G3488,G3487,G1440);
  nand GNAME3489(G3489,G7023,G1441);
  nand GNAME3490(G3490,G1347,G1442);
  nand GNAME3491(G3491,G1348,G1435);
  nand GNAME3492(G3492,G3417,G1349);
  nand GNAME3493(G3493,G3414,G21500);
  nand GNAME3494(G3494,G7026,G1444);
  nand GNAME3495(G3495,G25,G1446);
  nand GNAME3496(G3496,G9,G2275);
  nand GNAME3497(G3497,G3496,G3494,G3495);
  nand GNAME3498(G3498,G1447,G21426);
  nand GNAME3499(G3499,G3498,G2317);
  nand GNAME3500(G3500,G1443,G3499);
  nand GNAME3501(G3501,G3500,G1531);
  or GNAME3502(G3502,G2298,G1445);
  nand GNAME3503(G3503,G21426,G2275);
  nand GNAME3504(G3504,G3502,G3503);
  nand GNAME3505(G3505,G3497,G1448);
  nand GNAME3506(G3506,G7026,G1449);
  nand GNAME3507(G3507,G1325,G1450);
  nand GNAME3508(G3508,G1327,G2267);
  nand GNAME3509(G3509,G3504,G1328);
  nand GNAME3510(G3510,G3501,G21501);
  nand GNAME3511(G3511,G7029,G1444);
  nand GNAME3512(G3512,G26,G1446);
  nand GNAME3513(G3513,G10,G2275);
  nand GNAME3514(G3514,G3513,G3511,G3512);
  nand GNAME3515(G3515,G3514,G1448);
  nand GNAME3516(G3516,G7029,G1449);
  nand GNAME3517(G3517,G1329,G1450);
  nand GNAME3518(G3518,G1330,G2267);
  nand GNAME3519(G3519,G3504,G1331);
  nand GNAME3520(G3520,G3501,G21502);
  nand GNAME3521(G3521,G7032,G1444);
  nand GNAME3522(G3522,G27,G1446);
  nand GNAME3523(G3523,G11,G2275);
  nand GNAME3524(G3524,G3523,G3521,G3522);
  nand GNAME3525(G3525,G3524,G1448);
  nand GNAME3526(G3526,G7032,G1449);
  nand GNAME3527(G3527,G1332,G1450);
  nand GNAME3528(G3528,G1333,G2267);
  nand GNAME3529(G3529,G3504,G1334);
  nand GNAME3530(G3530,G3501,G21503);
  nand GNAME3531(G3531,G7035,G1444);
  nand GNAME3532(G3532,G28,G1446);
  nand GNAME3533(G3533,G12,G2275);
  nand GNAME3534(G3534,G3533,G3531,G3532);
  nand GNAME3535(G3535,G3534,G1448);
  nand GNAME3536(G3536,G7035,G1449);
  nand GNAME3537(G3537,G1335,G1450);
  nand GNAME3538(G3538,G1336,G2267);
  nand GNAME3539(G3539,G3504,G1337);
  nand GNAME3540(G3540,G3501,G21504);
  nand GNAME3541(G3541,G7038,G1444);
  nand GNAME3542(G3542,G29,G1446);
  nand GNAME3543(G3543,G13,G2275);
  nand GNAME3544(G3544,G3543,G3541,G3542);
  nand GNAME3545(G3545,G3544,G1448);
  nand GNAME3546(G3546,G7038,G1449);
  nand GNAME3547(G3547,G1338,G1450);
  nand GNAME3548(G3548,G1339,G2267);
  nand GNAME3549(G3549,G3504,G1340);
  nand GNAME3550(G3550,G3501,G21505);
  nand GNAME3551(G3551,G7041,G1444);
  nand GNAME3552(G3552,G30,G1446);
  nand GNAME3553(G3553,G14,G2275);
  nand GNAME3554(G3554,G3553,G3551,G3552);
  nand GNAME3555(G3555,G3554,G1448);
  nand GNAME3556(G3556,G7041,G1449);
  nand GNAME3557(G3557,G1341,G1450);
  nand GNAME3558(G3558,G1342,G2267);
  nand GNAME3559(G3559,G3504,G1343);
  nand GNAME3560(G3560,G3501,G21506);
  nand GNAME3561(G3561,G7044,G1444);
  nand GNAME3562(G3562,G31,G1446);
  nand GNAME3563(G3563,G15,G2275);
  nand GNAME3564(G3564,G3563,G3561,G3562);
  nand GNAME3565(G3565,G3564,G1448);
  nand GNAME3566(G3566,G7044,G1449);
  nand GNAME3567(G3567,G1344,G1450);
  nand GNAME3568(G3568,G1345,G2267);
  nand GNAME3569(G3569,G3504,G1346);
  nand GNAME3570(G3570,G3501,G21507);
  nand GNAME3571(G3571,G7047,G1444);
  nand GNAME3572(G3572,G32,G1446);
  nand GNAME3573(G3573,G16,G2275);
  nand GNAME3574(G3574,G3573,G3571,G3572);
  nand GNAME3575(G3575,G3574,G1448);
  nand GNAME3576(G3576,G7047,G1449);
  nand GNAME3577(G3577,G1347,G1450);
  nand GNAME3578(G3578,G1348,G2267);
  nand GNAME3579(G3579,G3504,G1349);
  nand GNAME3580(G3580,G3501,G21508);
  nand GNAME3581(G3581,G7050,G1453);
  nand GNAME3582(G3582,G25,G1455);
  nand GNAME3583(G3583,G9,G2274);
  nand GNAME3584(G3584,G3583,G3581,G3582);
  nand GNAME3585(G3585,G1456,G21426);
  nand GNAME3586(G3586,G3585,G2317);
  nand GNAME3587(G3587,G1452,G3586);
  nand GNAME3588(G3588,G3587,G1531);
  or GNAME3589(G3589,G2298,G1454);
  nand GNAME3590(G3590,G21426,G2274);
  nand GNAME3591(G3591,G3589,G3590);
  nand GNAME3592(G3592,G3584,G1457);
  nand GNAME3593(G3593,G7050,G1458);
  nand GNAME3594(G3594,G1325,G1459);
  nand GNAME3595(G3595,G1327,G2266);
  nand GNAME3596(G3596,G3591,G1328);
  nand GNAME3597(G3597,G3588,G21509);
  nand GNAME3598(G3598,G7053,G1453);
  nand GNAME3599(G3599,G26,G1455);
  nand GNAME3600(G3600,G10,G2274);
  nand GNAME3601(G3601,G3600,G3598,G3599);
  nand GNAME3602(G3602,G3601,G1457);
  nand GNAME3603(G3603,G7053,G1458);
  nand GNAME3604(G3604,G1329,G1459);
  nand GNAME3605(G3605,G1330,G2266);
  nand GNAME3606(G3606,G3591,G1331);
  nand GNAME3607(G3607,G3588,G21510);
  nand GNAME3608(G3608,G7056,G1453);
  nand GNAME3609(G3609,G27,G1455);
  nand GNAME3610(G3610,G11,G2274);
  nand GNAME3611(G3611,G3610,G3608,G3609);
  nand GNAME3612(G3612,G3611,G1457);
  nand GNAME3613(G3613,G7056,G1458);
  nand GNAME3614(G3614,G1332,G1459);
  nand GNAME3615(G3615,G1333,G2266);
  nand GNAME3616(G3616,G3591,G1334);
  nand GNAME3617(G3617,G3588,G21511);
  nand GNAME3618(G3618,G7059,G1453);
  nand GNAME3619(G3619,G28,G1455);
  nand GNAME3620(G3620,G12,G2274);
  nand GNAME3621(G3621,G3620,G3618,G3619);
  nand GNAME3622(G3622,G3621,G1457);
  nand GNAME3623(G3623,G7059,G1458);
  nand GNAME3624(G3624,G1335,G1459);
  nand GNAME3625(G3625,G1336,G2266);
  nand GNAME3626(G3626,G3591,G1337);
  nand GNAME3627(G3627,G3588,G21512);
  nand GNAME3628(G3628,G7062,G1453);
  nand GNAME3629(G3629,G29,G1455);
  nand GNAME3630(G3630,G13,G2274);
  nand GNAME3631(G3631,G3630,G3628,G3629);
  nand GNAME3632(G3632,G3631,G1457);
  nand GNAME3633(G3633,G7062,G1458);
  nand GNAME3634(G3634,G1338,G1459);
  nand GNAME3635(G3635,G1339,G2266);
  nand GNAME3636(G3636,G3591,G1340);
  nand GNAME3637(G3637,G3588,G21513);
  nand GNAME3638(G3638,G7065,G1453);
  nand GNAME3639(G3639,G30,G1455);
  nand GNAME3640(G3640,G14,G2274);
  nand GNAME3641(G3641,G3640,G3638,G3639);
  nand GNAME3642(G3642,G3641,G1457);
  nand GNAME3643(G3643,G7065,G1458);
  nand GNAME3644(G3644,G1341,G1459);
  nand GNAME3645(G3645,G1342,G2266);
  nand GNAME3646(G3646,G3591,G1343);
  nand GNAME3647(G3647,G3588,G21514);
  nand GNAME3648(G3648,G7068,G1453);
  nand GNAME3649(G3649,G31,G1455);
  nand GNAME3650(G3650,G15,G2274);
  nand GNAME3651(G3651,G3650,G3648,G3649);
  nand GNAME3652(G3652,G3651,G1457);
  nand GNAME3653(G3653,G7068,G1458);
  nand GNAME3654(G3654,G1344,G1459);
  nand GNAME3655(G3655,G1345,G2266);
  nand GNAME3656(G3656,G3591,G1346);
  nand GNAME3657(G3657,G3588,G21515);
  nand GNAME3658(G3658,G7071,G1453);
  nand GNAME3659(G3659,G32,G1455);
  nand GNAME3660(G3660,G16,G2274);
  nand GNAME3661(G3661,G3660,G3658,G3659);
  nand GNAME3662(G3662,G3661,G1457);
  nand GNAME3663(G3663,G7071,G1458);
  nand GNAME3664(G3664,G1347,G1459);
  nand GNAME3665(G3665,G1348,G2266);
  nand GNAME3666(G3666,G3591,G1349);
  nand GNAME3667(G3667,G3588,G21516);
  nand GNAME3668(G3668,G7074,G1461);
  nand GNAME3669(G3669,G25,G1463);
  nand GNAME3670(G3670,G9,G2273);
  nand GNAME3671(G3671,G3670,G3668,G3669);
  nand GNAME3672(G3672,G1464,G21426);
  nand GNAME3673(G3673,G3672,G2317);
  nand GNAME3674(G3674,G1460,G3673);
  nand GNAME3675(G3675,G3674,G1531);
  or GNAME3676(G3676,G2298,G1462);
  nand GNAME3677(G3677,G21426,G2273);
  nand GNAME3678(G3678,G3676,G3677);
  nand GNAME3679(G3679,G3671,G1465);
  nand GNAME3680(G3680,G7074,G1466);
  nand GNAME3681(G3681,G1325,G1467);
  nand GNAME3682(G3682,G1327,G2265);
  nand GNAME3683(G3683,G3678,G1328);
  nand GNAME3684(G3684,G3675,G21517);
  nand GNAME3685(G3685,G7077,G1461);
  nand GNAME3686(G3686,G26,G1463);
  nand GNAME3687(G3687,G10,G2273);
  nand GNAME3688(G3688,G3687,G3685,G3686);
  nand GNAME3689(G3689,G3688,G1465);
  nand GNAME3690(G3690,G7077,G1466);
  nand GNAME3691(G3691,G1329,G1467);
  nand GNAME3692(G3692,G1330,G2265);
  nand GNAME3693(G3693,G3678,G1331);
  nand GNAME3694(G3694,G3675,G21518);
  nand GNAME3695(G3695,G7080,G1461);
  nand GNAME3696(G3696,G27,G1463);
  nand GNAME3697(G3697,G11,G2273);
  nand GNAME3698(G3698,G3697,G3695,G3696);
  nand GNAME3699(G3699,G3698,G1465);
  nand GNAME3700(G3700,G7080,G1466);
  nand GNAME3701(G3701,G1332,G1467);
  nand GNAME3702(G3702,G1333,G2265);
  nand GNAME3703(G3703,G3678,G1334);
  nand GNAME3704(G3704,G3675,G21519);
  nand GNAME3705(G3705,G7083,G1461);
  nand GNAME3706(G3706,G28,G1463);
  nand GNAME3707(G3707,G12,G2273);
  nand GNAME3708(G3708,G3707,G3705,G3706);
  nand GNAME3709(G3709,G3708,G1465);
  nand GNAME3710(G3710,G7083,G1466);
  nand GNAME3711(G3711,G1335,G1467);
  nand GNAME3712(G3712,G1336,G2265);
  nand GNAME3713(G3713,G3678,G1337);
  nand GNAME3714(G3714,G3675,G21520);
  nand GNAME3715(G3715,G7086,G1461);
  nand GNAME3716(G3716,G29,G1463);
  nand GNAME3717(G3717,G13,G2273);
  nand GNAME3718(G3718,G3717,G3715,G3716);
  nand GNAME3719(G3719,G3718,G1465);
  nand GNAME3720(G3720,G7086,G1466);
  nand GNAME3721(G3721,G1338,G1467);
  nand GNAME3722(G3722,G1339,G2265);
  nand GNAME3723(G3723,G3678,G1340);
  nand GNAME3724(G3724,G3675,G21521);
  nand GNAME3725(G3725,G7089,G1461);
  nand GNAME3726(G3726,G30,G1463);
  nand GNAME3727(G3727,G14,G2273);
  nand GNAME3728(G3728,G3727,G3725,G3726);
  nand GNAME3729(G3729,G3728,G1465);
  nand GNAME3730(G3730,G7089,G1466);
  nand GNAME3731(G3731,G1341,G1467);
  nand GNAME3732(G3732,G1342,G2265);
  nand GNAME3733(G3733,G3678,G1343);
  nand GNAME3734(G3734,G3675,G21522);
  nand GNAME3735(G3735,G7092,G1461);
  nand GNAME3736(G3736,G31,G1463);
  nand GNAME3737(G3737,G15,G2273);
  nand GNAME3738(G3738,G3737,G3735,G3736);
  nand GNAME3739(G3739,G3738,G1465);
  nand GNAME3740(G3740,G7092,G1466);
  nand GNAME3741(G3741,G1344,G1467);
  nand GNAME3742(G3742,G1345,G2265);
  nand GNAME3743(G3743,G3678,G1346);
  nand GNAME3744(G3744,G3675,G21523);
  nand GNAME3745(G3745,G7095,G1461);
  nand GNAME3746(G3746,G32,G1463);
  nand GNAME3747(G3747,G16,G2273);
  nand GNAME3748(G3748,G3747,G3745,G3746);
  nand GNAME3749(G3749,G3748,G1465);
  nand GNAME3750(G3750,G7095,G1466);
  nand GNAME3751(G3751,G1347,G1467);
  nand GNAME3752(G3752,G1348,G2265);
  nand GNAME3753(G3753,G3678,G1349);
  nand GNAME3754(G3754,G3675,G21524);
  nand GNAME3755(G3755,G7098,G1470);
  nand GNAME3756(G3756,G25,G1472);
  nand GNAME3757(G3757,G9,G2272);
  nand GNAME3758(G3758,G3757,G3755,G3756);
  nand GNAME3759(G3759,G1473,G21426);
  nand GNAME3760(G3760,G3759,G2317);
  nand GNAME3761(G3761,G1469,G3760);
  nand GNAME3762(G3762,G3761,G1531);
  or GNAME3763(G3763,G2298,G1471);
  nand GNAME3764(G3764,G21426,G2272);
  nand GNAME3765(G3765,G3763,G3764);
  nand GNAME3766(G3766,G3758,G1474);
  nand GNAME3767(G3767,G7098,G1475);
  nand GNAME3768(G3768,G1325,G1476);
  nand GNAME3769(G3769,G1327,G2264);
  nand GNAME3770(G3770,G3765,G1328);
  nand GNAME3771(G3771,G3762,G21525);
  nand GNAME3772(G3772,G7101,G1470);
  nand GNAME3773(G3773,G26,G1472);
  nand GNAME3774(G3774,G10,G2272);
  nand GNAME3775(G3775,G3774,G3772,G3773);
  nand GNAME3776(G3776,G3775,G1474);
  nand GNAME3777(G3777,G7101,G1475);
  nand GNAME3778(G3778,G1329,G1476);
  nand GNAME3779(G3779,G1330,G2264);
  nand GNAME3780(G3780,G3765,G1331);
  nand GNAME3781(G3781,G3762,G21526);
  nand GNAME3782(G3782,G7104,G1470);
  nand GNAME3783(G3783,G27,G1472);
  nand GNAME3784(G3784,G11,G2272);
  nand GNAME3785(G3785,G3784,G3782,G3783);
  nand GNAME3786(G3786,G3785,G1474);
  nand GNAME3787(G3787,G7104,G1475);
  nand GNAME3788(G3788,G1332,G1476);
  nand GNAME3789(G3789,G1333,G2264);
  nand GNAME3790(G3790,G3765,G1334);
  nand GNAME3791(G3791,G3762,G21527);
  nand GNAME3792(G3792,G7107,G1470);
  nand GNAME3793(G3793,G28,G1472);
  nand GNAME3794(G3794,G12,G2272);
  nand GNAME3795(G3795,G3794,G3792,G3793);
  nand GNAME3796(G3796,G3795,G1474);
  nand GNAME3797(G3797,G7107,G1475);
  nand GNAME3798(G3798,G1335,G1476);
  nand GNAME3799(G3799,G1336,G2264);
  nand GNAME3800(G3800,G3765,G1337);
  nand GNAME3801(G3801,G3762,G21528);
  nand GNAME3802(G3802,G7110,G1470);
  nand GNAME3803(G3803,G29,G1472);
  nand GNAME3804(G3804,G13,G2272);
  nand GNAME3805(G3805,G3804,G3802,G3803);
  nand GNAME3806(G3806,G3805,G1474);
  nand GNAME3807(G3807,G7110,G1475);
  nand GNAME3808(G3808,G1338,G1476);
  nand GNAME3809(G3809,G1339,G2264);
  nand GNAME3810(G3810,G3765,G1340);
  nand GNAME3811(G3811,G3762,G21529);
  nand GNAME3812(G3812,G7113,G1470);
  nand GNAME3813(G3813,G30,G1472);
  nand GNAME3814(G3814,G14,G2272);
  nand GNAME3815(G3815,G3814,G3812,G3813);
  nand GNAME3816(G3816,G3815,G1474);
  nand GNAME3817(G3817,G7113,G1475);
  nand GNAME3818(G3818,G1341,G1476);
  nand GNAME3819(G3819,G1342,G2264);
  nand GNAME3820(G3820,G3765,G1343);
  nand GNAME3821(G3821,G3762,G21530);
  nand GNAME3822(G3822,G7116,G1470);
  nand GNAME3823(G3823,G31,G1472);
  nand GNAME3824(G3824,G15,G2272);
  nand GNAME3825(G3825,G3824,G3822,G3823);
  nand GNAME3826(G3826,G3825,G1474);
  nand GNAME3827(G3827,G7116,G1475);
  nand GNAME3828(G3828,G1344,G1476);
  nand GNAME3829(G3829,G1345,G2264);
  nand GNAME3830(G3830,G3765,G1346);
  nand GNAME3831(G3831,G3762,G21531);
  nand GNAME3832(G3832,G7119,G1470);
  nand GNAME3833(G3833,G32,G1472);
  nand GNAME3834(G3834,G16,G2272);
  nand GNAME3835(G3835,G3834,G3832,G3833);
  nand GNAME3836(G3836,G3835,G1474);
  nand GNAME3837(G3837,G7119,G1475);
  nand GNAME3838(G3838,G1347,G1476);
  nand GNAME3839(G3839,G1348,G2264);
  nand GNAME3840(G3840,G3765,G1349);
  nand GNAME3841(G3841,G3762,G21532);
  nand GNAME3842(G3842,G7122,G1478);
  nand GNAME3843(G3843,G25,G1480);
  nand GNAME3844(G3844,G9,G2271);
  nand GNAME3845(G3845,G3844,G3842,G3843);
  nand GNAME3846(G3846,G1481,G21426);
  nand GNAME3847(G3847,G3846,G2317);
  nand GNAME3848(G3848,G1477,G3847);
  nand GNAME3849(G3849,G3848,G1531);
  or GNAME3850(G3850,G2298,G1479);
  nand GNAME3851(G3851,G21426,G2271);
  nand GNAME3852(G3852,G3850,G3851);
  nand GNAME3853(G3853,G3845,G1482);
  nand GNAME3854(G3854,G7122,G1483);
  nand GNAME3855(G3855,G1325,G1484);
  nand GNAME3856(G3856,G1327,G2263);
  nand GNAME3857(G3857,G3852,G1328);
  nand GNAME3858(G3858,G3849,G21533);
  nand GNAME3859(G3859,G7125,G1478);
  nand GNAME3860(G3860,G26,G1480);
  nand GNAME3861(G3861,G10,G2271);
  nand GNAME3862(G3862,G3861,G3859,G3860);
  nand GNAME3863(G3863,G3862,G1482);
  nand GNAME3864(G3864,G7125,G1483);
  nand GNAME3865(G3865,G1329,G1484);
  nand GNAME3866(G3866,G1330,G2263);
  nand GNAME3867(G3867,G3852,G1331);
  nand GNAME3868(G3868,G3849,G21534);
  nand GNAME3869(G3869,G7128,G1478);
  nand GNAME3870(G3870,G27,G1480);
  nand GNAME3871(G3871,G11,G2271);
  nand GNAME3872(G3872,G3871,G3869,G3870);
  nand GNAME3873(G3873,G3872,G1482);
  nand GNAME3874(G3874,G7128,G1483);
  nand GNAME3875(G3875,G1332,G1484);
  nand GNAME3876(G3876,G1333,G2263);
  nand GNAME3877(G3877,G3852,G1334);
  nand GNAME3878(G3878,G3849,G21535);
  nand GNAME3879(G3879,G7131,G1478);
  nand GNAME3880(G3880,G28,G1480);
  nand GNAME3881(G3881,G12,G2271);
  nand GNAME3882(G3882,G3881,G3879,G3880);
  nand GNAME3883(G3883,G3882,G1482);
  nand GNAME3884(G3884,G7131,G1483);
  nand GNAME3885(G3885,G1335,G1484);
  nand GNAME3886(G3886,G1336,G2263);
  nand GNAME3887(G3887,G3852,G1337);
  nand GNAME3888(G3888,G3849,G21536);
  nand GNAME3889(G3889,G7134,G1478);
  nand GNAME3890(G3890,G29,G1480);
  nand GNAME3891(G3891,G13,G2271);
  nand GNAME3892(G3892,G3891,G3889,G3890);
  nand GNAME3893(G3893,G3892,G1482);
  nand GNAME3894(G3894,G7134,G1483);
  nand GNAME3895(G3895,G1338,G1484);
  nand GNAME3896(G3896,G1339,G2263);
  nand GNAME3897(G3897,G3852,G1340);
  nand GNAME3898(G3898,G3849,G21537);
  nand GNAME3899(G3899,G7137,G1478);
  nand GNAME3900(G3900,G30,G1480);
  nand GNAME3901(G3901,G14,G2271);
  nand GNAME3902(G3902,G3901,G3899,G3900);
  nand GNAME3903(G3903,G3902,G1482);
  nand GNAME3904(G3904,G7137,G1483);
  nand GNAME3905(G3905,G1341,G1484);
  nand GNAME3906(G3906,G1342,G2263);
  nand GNAME3907(G3907,G3852,G1343);
  nand GNAME3908(G3908,G3849,G21538);
  nand GNAME3909(G3909,G7140,G1478);
  nand GNAME3910(G3910,G31,G1480);
  nand GNAME3911(G3911,G15,G2271);
  nand GNAME3912(G3912,G3911,G3909,G3910);
  nand GNAME3913(G3913,G3912,G1482);
  nand GNAME3914(G3914,G7140,G1483);
  nand GNAME3915(G3915,G1344,G1484);
  nand GNAME3916(G3916,G1345,G2263);
  nand GNAME3917(G3917,G3852,G1346);
  nand GNAME3918(G3918,G3849,G21539);
  nand GNAME3919(G3919,G7143,G1478);
  nand GNAME3920(G3920,G32,G1480);
  nand GNAME3921(G3921,G16,G2271);
  nand GNAME3922(G3922,G3921,G3919,G3920);
  nand GNAME3923(G3923,G3922,G1482);
  nand GNAME3924(G3924,G7143,G1483);
  nand GNAME3925(G3925,G1347,G1484);
  nand GNAME3926(G3926,G1348,G2263);
  nand GNAME3927(G3927,G3852,G1349);
  nand GNAME3928(G3928,G3849,G21540);
  nand GNAME3929(G3929,G7146,G1486);
  nand GNAME3930(G3930,G25,G1488);
  nand GNAME3931(G3931,G9,G2270);
  nand GNAME3932(G3932,G3931,G3929,G3930);
  nand GNAME3933(G3933,G1489,G21426);
  nand GNAME3934(G3934,G3933,G2317);
  nand GNAME3935(G3935,G1485,G3934);
  nand GNAME3936(G3936,G3935,G1531);
  or GNAME3937(G3937,G2298,G1487);
  nand GNAME3938(G3938,G21426,G2270);
  nand GNAME3939(G3939,G3937,G3938);
  nand GNAME3940(G3940,G3932,G1490);
  nand GNAME3941(G3941,G7146,G1491);
  nand GNAME3942(G3942,G1325,G1492);
  nand GNAME3943(G3943,G1327,G2262);
  nand GNAME3944(G3944,G3939,G1328);
  nand GNAME3945(G3945,G3936,G21541);
  nand GNAME3946(G3946,G7149,G1486);
  nand GNAME3947(G3947,G26,G1488);
  nand GNAME3948(G3948,G10,G2270);
  nand GNAME3949(G3949,G3948,G3946,G3947);
  nand GNAME3950(G3950,G3949,G1490);
  nand GNAME3951(G3951,G7149,G1491);
  nand GNAME3952(G3952,G1329,G1492);
  nand GNAME3953(G3953,G1330,G2262);
  nand GNAME3954(G3954,G3939,G1331);
  nand GNAME3955(G3955,G3936,G21542);
  nand GNAME3956(G3956,G7152,G1486);
  nand GNAME3957(G3957,G27,G1488);
  nand GNAME3958(G3958,G11,G2270);
  nand GNAME3959(G3959,G3958,G3956,G3957);
  nand GNAME3960(G3960,G3959,G1490);
  nand GNAME3961(G3961,G7152,G1491);
  nand GNAME3962(G3962,G1332,G1492);
  nand GNAME3963(G3963,G1333,G2262);
  nand GNAME3964(G3964,G3939,G1334);
  nand GNAME3965(G3965,G3936,G21543);
  nand GNAME3966(G3966,G7155,G1486);
  nand GNAME3967(G3967,G28,G1488);
  nand GNAME3968(G3968,G12,G2270);
  nand GNAME3969(G3969,G3968,G3966,G3967);
  nand GNAME3970(G3970,G3969,G1490);
  nand GNAME3971(G3971,G7155,G1491);
  nand GNAME3972(G3972,G1335,G1492);
  nand GNAME3973(G3973,G1336,G2262);
  nand GNAME3974(G3974,G3939,G1337);
  nand GNAME3975(G3975,G3936,G21544);
  nand GNAME3976(G3976,G7158,G1486);
  nand GNAME3977(G3977,G29,G1488);
  nand GNAME3978(G3978,G13,G2270);
  nand GNAME3979(G3979,G3978,G3976,G3977);
  nand GNAME3980(G3980,G3979,G1490);
  nand GNAME3981(G3981,G7158,G1491);
  nand GNAME3982(G3982,G1338,G1492);
  nand GNAME3983(G3983,G1339,G2262);
  nand GNAME3984(G3984,G3939,G1340);
  nand GNAME3985(G3985,G3936,G21545);
  nand GNAME3986(G3986,G7161,G1486);
  nand GNAME3987(G3987,G30,G1488);
  nand GNAME3988(G3988,G14,G2270);
  nand GNAME3989(G3989,G3988,G3986,G3987);
  nand GNAME3990(G3990,G3989,G1490);
  nand GNAME3991(G3991,G7161,G1491);
  nand GNAME3992(G3992,G1341,G1492);
  nand GNAME3993(G3993,G1342,G2262);
  nand GNAME3994(G3994,G3939,G1343);
  nand GNAME3995(G3995,G3936,G21546);
  nand GNAME3996(G3996,G7164,G1486);
  nand GNAME3997(G3997,G31,G1488);
  nand GNAME3998(G3998,G15,G2270);
  nand GNAME3999(G3999,G3998,G3996,G3997);
  nand GNAME4000(G4000,G3999,G1490);
  nand GNAME4001(G4001,G7164,G1491);
  nand GNAME4002(G4002,G1344,G1492);
  nand GNAME4003(G4003,G1345,G2262);
  nand GNAME4004(G4004,G3939,G1346);
  nand GNAME4005(G4005,G3936,G21547);
  nand GNAME4006(G4006,G7167,G1486);
  nand GNAME4007(G4007,G32,G1488);
  nand GNAME4008(G4008,G16,G2270);
  nand GNAME4009(G4009,G4008,G4006,G4007);
  nand GNAME4010(G4010,G4009,G1490);
  nand GNAME4011(G4011,G7167,G1491);
  nand GNAME4012(G4012,G1347,G1492);
  nand GNAME4013(G4013,G1348,G2262);
  nand GNAME4014(G4014,G3939,G1349);
  nand GNAME4015(G4015,G3936,G21548);
  nand GNAME4016(G4016,G7170,G1494);
  nand GNAME4017(G4017,G25,G1496);
  nand GNAME4018(G4018,G9,G2269);
  nand GNAME4019(G4019,G4018,G4016,G4017);
  nand GNAME4020(G4020,G1497,G21426);
  nand GNAME4021(G4021,G4020,G2317);
  nand GNAME4022(G4022,G1493,G4021);
  nand GNAME4023(G4023,G4022,G1531);
  or GNAME4024(G4024,G2298,G1495);
  nand GNAME4025(G4025,G21426,G2269);
  nand GNAME4026(G4026,G4024,G4025);
  nand GNAME4027(G4027,G4019,G1498);
  nand GNAME4028(G4028,G7170,G1499);
  nand GNAME4029(G4029,G1325,G1500);
  nand GNAME4030(G4030,G1327,G2261);
  nand GNAME4031(G4031,G4026,G1328);
  nand GNAME4032(G4032,G4023,G21549);
  nand GNAME4033(G4033,G7173,G1494);
  nand GNAME4034(G4034,G26,G1496);
  nand GNAME4035(G4035,G10,G2269);
  nand GNAME4036(G4036,G4035,G4033,G4034);
  nand GNAME4037(G4037,G4036,G1498);
  nand GNAME4038(G4038,G7173,G1499);
  nand GNAME4039(G4039,G1329,G1500);
  nand GNAME4040(G4040,G1330,G2261);
  nand GNAME4041(G4041,G4026,G1331);
  nand GNAME4042(G4042,G4023,G21550);
  nand GNAME4043(G4043,G7176,G1494);
  nand GNAME4044(G4044,G27,G1496);
  nand GNAME4045(G4045,G11,G2269);
  nand GNAME4046(G4046,G4045,G4043,G4044);
  nand GNAME4047(G4047,G4046,G1498);
  nand GNAME4048(G4048,G7176,G1499);
  nand GNAME4049(G4049,G1332,G1500);
  nand GNAME4050(G4050,G1333,G2261);
  nand GNAME4051(G4051,G4026,G1334);
  nand GNAME4052(G4052,G4023,G21551);
  nand GNAME4053(G4053,G7179,G1494);
  nand GNAME4054(G4054,G28,G1496);
  nand GNAME4055(G4055,G12,G2269);
  nand GNAME4056(G4056,G4055,G4053,G4054);
  nand GNAME4057(G4057,G4056,G1498);
  nand GNAME4058(G4058,G7179,G1499);
  nand GNAME4059(G4059,G1335,G1500);
  nand GNAME4060(G4060,G1336,G2261);
  nand GNAME4061(G4061,G4026,G1337);
  nand GNAME4062(G4062,G4023,G21552);
  nand GNAME4063(G4063,G7182,G1494);
  nand GNAME4064(G4064,G29,G1496);
  nand GNAME4065(G4065,G13,G2269);
  nand GNAME4066(G4066,G4065,G4063,G4064);
  nand GNAME4067(G4067,G4066,G1498);
  nand GNAME4068(G4068,G7182,G1499);
  nand GNAME4069(G4069,G1338,G1500);
  nand GNAME4070(G4070,G1339,G2261);
  nand GNAME4071(G4071,G4026,G1340);
  nand GNAME4072(G4072,G4023,G21553);
  nand GNAME4073(G4073,G7185,G1494);
  nand GNAME4074(G4074,G30,G1496);
  nand GNAME4075(G4075,G14,G2269);
  nand GNAME4076(G4076,G4075,G4073,G4074);
  nand GNAME4077(G4077,G4076,G1498);
  nand GNAME4078(G4078,G7185,G1499);
  nand GNAME4079(G4079,G1341,G1500);
  nand GNAME4080(G4080,G1342,G2261);
  nand GNAME4081(G4081,G4026,G1343);
  nand GNAME4082(G4082,G4023,G21554);
  nand GNAME4083(G4083,G7188,G1494);
  nand GNAME4084(G4084,G31,G1496);
  nand GNAME4085(G4085,G15,G2269);
  nand GNAME4086(G4086,G4085,G4083,G4084);
  nand GNAME4087(G4087,G4086,G1498);
  nand GNAME4088(G4088,G7188,G1499);
  nand GNAME4089(G4089,G1344,G1500);
  nand GNAME4090(G4090,G1345,G2261);
  nand GNAME4091(G4091,G4026,G1346);
  nand GNAME4092(G4092,G4023,G21555);
  nand GNAME4093(G4093,G7191,G1494);
  nand GNAME4094(G4094,G32,G1496);
  nand GNAME4095(G4095,G16,G2269);
  nand GNAME4096(G4096,G4095,G4093,G4094);
  nand GNAME4097(G4097,G4096,G1498);
  nand GNAME4098(G4098,G7191,G1499);
  nand GNAME4099(G4099,G1347,G1500);
  nand GNAME4100(G4100,G1348,G2261);
  nand GNAME4101(G4101,G4026,G1349);
  nand GNAME4102(G4102,G4023,G21556);
  nand GNAME4103(G4103,G2600,G2477);
  nand GNAME4104(G4104,G1192,G2545);
  nand GNAME4105(G4105,G4104,G1501);
  nand GNAME4106(G4106,G1556,G1247);
  nand GNAME4107(G4107,G1255,G4106,G2460);
  nand GNAME4108(G4108,G1202,G2325);
  nand GNAME4109(G4109,G2609,G4107,G4108);
  or GNAME4110(G4110,G1502,G35,G1190);
  nand GNAME4111(G4111,G4109,G7326);
  nand GNAME4112(G4112,G2257,G1506);
  nand GNAME4113(G4113,G2340,G1233);
  nand GNAME4114(G4114,G1212,G2340);
  nand GNAME4115(G4115,G4114,G21558);
  nand GNAME4116(G4116,G1215,G7207,G7208);
  nand GNAME4117(G4117,G4116,G7207);
  not GNAME4118(G4118,G1518);
  nand GNAME4119(G4119,G1244,G1514);
  nand GNAME4120(G4120,G4119,G1515);
  nand GNAME4121(G4121,G1192,G4120);
  nand GNAME4122(G4122,G1563,G1504,G2326,G4121);
  nand GNAME4123(G4123,G1249,G1516);
  or GNAME4124(G4124,G2477,G1517);
  nand GNAME4125(G4125,G2545,G1262);
  nand GNAME4126(G4126,G1249,G1240);
  nand GNAME4127(G4127,G2608,G1250);
  nand GNAME4128(G4128,G2311,G1518);
  nand GNAME4129(G4129,G6750,G7198,G7199);
  and GNAME4130(G4130,G4118,G1509);
  or GNAME4131(G4131,G4130,G1260);
  nand GNAME4132(G4132,G1238,G1266);
  nand GNAME4133(G4133,G4132,G1522);
  nand GNAME4134(G4134,G2321,G1190,G1717);
  nand GNAME4135(G4135,G1556,G1572);
  nand GNAME4136(G4136,G4135,G1729);
  nand GNAME4137(G4137,G4134,G6804);
  nand GNAME4138(G4138,G4133,G7443);
  nand GNAME4139(G4139,G4122,G7779);
  nand GNAME4140(G4140,G1523,G1524);
  nand GNAME4141(G4141,G7204,G1525);
  nand GNAME4142(G4142,G1934,G4138,G4136,G4139);
  nand GNAME4143(G4143,G1507,G7779);
  nand GNAME4144(G4144,G4142,G1283);
  nand GNAME4145(G4145,G4143,G4144);
  nand GNAME4146(G4146,G2348,G7209);
  nand GNAME4147(G4147,G4135,G1739);
  nand GNAME4148(G4148,G4134,G2259);
  nand GNAME4149(G4149,G4133,G7440);
  nand GNAME4150(G4150,G4122,G7776);
  nand GNAME4151(G4151,G1523,G1730);
  nand GNAME4152(G4152,G1525,G2260);
  nand GNAME4153(G4153,G1935,G4149,G4147,G4150);
  nand GNAME4154(G4154,G2259,G1526);
  nand GNAME4155(G4155,G1507,G7776);
  nand GNAME4156(G4156,G4153,G1283);
  nand GNAME4157(G4157,G4156,G4154,G4155);
  not GNAME4158(G4158,G1688);
  nand GNAME4159(G4159,G21561,G2511);
  not GNAME4160(G4160,G1193);
  or GNAME4161(G4161,G1219,G4160);
  nand GNAME4162(G4162,G4161,G1523);
  nand GNAME4163(G4163,G4135,G1728);
  nand GNAME4164(G4164,G4134,G1727);
  nand GNAME4165(G4165,G4133,G7482);
  nand GNAME4166(G4166,G4122,G7824);
  nand GNAME4167(G4167,G1688,G1525);
  nand GNAME4168(G4168,G1936,G4164,G4166,G4163);
  nand GNAME4169(G4169,G1727,G1526);
  nand GNAME4170(G4170,G1507,G7824);
  nand GNAME4171(G4171,G4168,G1283);
  nand GNAME4172(G4172,G4171,G4169,G4170);
  nand GNAME4173(G4173,G1210,G1263);
  nand GNAME4174(G4174,G4135,G2277);
  nand GNAME4175(G4175,G4134,G2258);
  nand GNAME4176(G4176,G4133,G7467);
  nand GNAME4177(G4177,G4122,G7809);
  nand GNAME4178(G4178,G4176,G4177,G4175,G4173,G4174);
  nand GNAME4179(G4179,G1303,G6787);
  nand GNAME4180(G4180,G1507,G7809);
  nand GNAME4181(G4181,G4179,G21427);
  nand GNAME4182(G4182,G4178,G1283);
  nand GNAME4183(G4183,G4182,G4180,G4181);
  nand GNAME4184(G4184,G1282,G1274);
  nand GNAME4185(G4185,G1209,G2298);
  nand GNAME4186(G4186,G4185,G2306);
  nand GNAME4187(G4187,G6804,G1533);
  nand GNAME4188(G4188,G7443,G1534);
  or GNAME4189(G4189,G1287,G1532);
  nand GNAME4190(G4190,G2259,G1533);
  nand GNAME4191(G4191,G7440,G1534);
  or GNAME4192(G4192,G1286,G1532);
  nand GNAME4193(G4193,G1727,G1533);
  nand GNAME4194(G4194,G7482,G1534);
  or GNAME4195(G4195,G1284,G1532);
  nand GNAME4196(G4196,G1279,G2258);
  nand GNAME4197(G4197,G4186,G7467);
  nand GNAME4198(G4198,G21428,G7326);
  nand GNAME4199(G4199,G4198,G4196,G4197);
  nand GNAME4200(G4200,G2545,G2477);
  nand GNAME4201(G4201,G4200,G2596);
  nand GNAME4202(G4202,G1255,G1204,G4201);
  nand GNAME4203(G4203,G2494,G2346,G4202);
  nand GNAME4204(G4204,G2494,G1202,G1238);
  nand GNAME4205(G4205,G4204,G2528);
  nand GNAME4206(G4206,G8101,G4205,G2596);
  nand GNAME4207(G4207,G4203,G7326);
  nand GNAME4208(G4208,G1505,G4206,G4207);
  nand GNAME4209(G4209,G4208,G1506);
  nand GNAME4210(G4210,G1717,G2321,G1572,G1522);
  nand GNAME4211(G4211,G1504,G1937,G2327,G1556,G2326);
  nand GNAME4212(G4212,G2318,G1190,G1563,G7290);
  nand GNAME4213(G4213,G1537,G8258);
  nand GNAME4214(G4214,G7467,G1538);
  nand GNAME4215(G4215,G7809,G1539);
  nand GNAME4216(G4216,G1540,G8709);
  nand GNAME4217(G4217,G1541,G21758);
  nand GNAME4218(G4218,G21567,G1543);
  nand GNAME4219(G4219,G1537,G8273);
  nand GNAME4220(G4220,G7482,G1538);
  nand GNAME4221(G4221,G7824,G1539);
  nand GNAME4222(G4222,G1540,G8762);
  nand GNAME4223(G4223,G21759,G1541);
  nand GNAME4224(G4224,G1543,G21568);
  nand GNAME4225(G4225,G1537,G8208);
  nand GNAME4226(G4226,G7440,G1538);
  nand GNAME4227(G4227,G7776,G1539);
  nand GNAME4228(G4228,G1540,G8708);
  nand GNAME4229(G4229,G21760,G1541);
  nand GNAME4230(G4230,G1543,G21569);
  nand GNAME4231(G4231,G1537,G8211);
  nand GNAME4232(G4232,G7443,G1538);
  nand GNAME4233(G4233,G7779,G1539);
  nand GNAME4234(G4234,G1540,G8782);
  nand GNAME4235(G4235,G21761,G1541);
  nand GNAME4236(G4236,G1543,G21570);
  nand GNAME4237(G4237,G1537,G8262);
  nand GNAME4238(G4238,G1538,G7471);
  nand GNAME4239(G4239,G7813,G1539);
  nand GNAME4240(G4240,G1540,G8759);
  nand GNAME4241(G4241,G21762,G1541);
  nand GNAME4242(G4242,G1543,G21571);
  nand GNAME4243(G4243,G1537,G8261);
  nand GNAME4244(G4244,G1538,G7470);
  nand GNAME4245(G4245,G1539,G7812);
  nand GNAME4246(G4246,G1540,G8758);
  nand GNAME4247(G4247,G21763,G1541);
  nand GNAME4248(G4248,G1543,G21572);
  nand GNAME4249(G4249,G1537,G8212);
  nand GNAME4250(G4250,G1538,G7444);
  nand GNAME4251(G4251,G1539,G7780);
  nand GNAME4252(G4252,G1540,G8757);
  nand GNAME4253(G4253,G21764,G1541);
  nand GNAME4254(G4254,G1543,G21573);
  nand GNAME4255(G4255,G1537,G8213);
  nand GNAME4256(G4256,G1538,G7445);
  nand GNAME4257(G4257,G1539,G7781);
  nand GNAME4258(G4258,G1540,G8756);
  nand GNAME4259(G4259,G21765,G1541);
  nand GNAME4260(G4260,G1543,G21574);
  nand GNAME4261(G4261,G1537,G8260);
  nand GNAME4262(G4262,G1538,G7469);
  nand GNAME4263(G4263,G1539,G7811);
  nand GNAME4264(G4264,G1540,G8755);
  nand GNAME4265(G4265,G21766,G1541);
  nand GNAME4266(G4266,G1543,G21575);
  nand GNAME4267(G4267,G1537,G8259);
  nand GNAME4268(G4268,G1538,G7468);
  nand GNAME4269(G4269,G1539,G7810);
  nand GNAME4270(G4270,G1540,G8754);
  nand GNAME4271(G4271,G21767,G1541);
  nand GNAME4272(G4272,G1543,G21576);
  nand GNAME4273(G4273,G1537,G8205);
  nand GNAME4274(G4274,G1538,G7437);
  nand GNAME4275(G4275,G1539,G7773);
  nand GNAME4276(G4276,G1540,G8769);
  nand GNAME4277(G4277,G21768,G1541);
  nand GNAME4278(G4278,G1543,G21577);
  nand GNAME4279(G4279,G1537,G8206);
  nand GNAME4280(G4280,G1538,G7438);
  nand GNAME4281(G4281,G1539,G7774);
  nand GNAME4282(G4282,G1540,G8768);
  nand GNAME4283(G4283,G21769,G1541);
  nand GNAME4284(G4284,G1543,G21578);
  nand GNAME4285(G4285,G1537,G8280);
  nand GNAME4286(G4286,G1538,G7489);
  nand GNAME4287(G4287,G1539,G7831);
  nand GNAME4288(G4288,G1540,G8767);
  nand GNAME4289(G4289,G21770,G1541);
  nand GNAME4290(G4290,G1543,G21579);
  nand GNAME4291(G4291,G1537,G8279);
  nand GNAME4292(G4292,G1538,G7488);
  nand GNAME4293(G4293,G1539,G7830);
  nand GNAME4294(G4294,G1540,G8766);
  nand GNAME4295(G4295,G21771,G1541);
  nand GNAME4296(G4296,G1543,G21580);
  nand GNAME4297(G4297,G1537,G8207);
  nand GNAME4298(G4298,G1538,G7439);
  nand GNAME4299(G4299,G1539,G7775);
  nand GNAME4300(G4300,G1540,G8765);
  nand GNAME4301(G4301,G21772,G1541);
  nand GNAME4302(G4302,G1543,G21581);
  nand GNAME4303(G4303,G1537,G8278);
  nand GNAME4304(G4304,G1538,G7487);
  nand GNAME4305(G4305,G1539,G7829);
  nand GNAME4306(G4306,G1540,G8764);
  nand GNAME4307(G4307,G21773,G1541);
  nand GNAME4308(G4308,G1543,G21582);
  nand GNAME4309(G4309,G1537,G8277);
  nand GNAME4310(G4310,G1538,G7486);
  nand GNAME4311(G4311,G1539,G7828);
  nand GNAME4312(G4312,G1540,G8763);
  nand GNAME4313(G4313,G21774,G1541);
  nand GNAME4314(G4314,G1543,G21583);
  nand GNAME4315(G4315,G1537,G8276);
  nand GNAME4316(G4316,G1538,G7485);
  nand GNAME4317(G4317,G1539,G7827);
  nand GNAME4318(G4318,G1540,G8777);
  nand GNAME4319(G4319,G21775,G1541);
  nand GNAME4320(G4320,G1543,G21584);
  nand GNAME4321(G4321,G1537,G8275);
  nand GNAME4322(G4322,G1538,G7484);
  nand GNAME4323(G4323,G1539,G7826);
  nand GNAME4324(G4324,G1540,G8776);
  nand GNAME4325(G4325,G21776,G1541);
  nand GNAME4326(G4326,G1543,G21585);
  nand GNAME4327(G4327,G1537,G8274);
  nand GNAME4328(G4328,G1538,G7483);
  nand GNAME4329(G4329,G1539,G7825);
  nand GNAME4330(G4330,G1540,G8775);
  nand GNAME4331(G4331,G21777,G1541);
  nand GNAME4332(G4332,G1543,G21586);
  nand GNAME4333(G4333,G1537,G8272);
  nand GNAME4334(G4334,G1538,G7481);
  nand GNAME4335(G4335,G1539,G7823);
  nand GNAME4336(G4336,G1540,G8774);
  nand GNAME4337(G4337,G21778,G1541);
  nand GNAME4338(G4338,G1543,G21587);
  nand GNAME4339(G4339,G1537,G8271);
  nand GNAME4340(G4340,G1538,G7480);
  nand GNAME4341(G4341,G1539,G7822);
  nand GNAME4342(G4342,G1540,G8773);
  nand GNAME4343(G4343,G21779,G1541);
  nand GNAME4344(G4344,G1543,G21588);
  nand GNAME4345(G4345,G1537,G8270);
  nand GNAME4346(G4346,G1538,G7479);
  nand GNAME4347(G4347,G1539,G7821);
  nand GNAME4348(G4348,G1540,G8772);
  nand GNAME4349(G4349,G21780,G1541);
  nand GNAME4350(G4350,G1543,G21589);
  nand GNAME4351(G4351,G1537,G8269);
  nand GNAME4352(G4352,G1538,G7478);
  nand GNAME4353(G4353,G1539,G7820);
  nand GNAME4354(G4354,G1540,G8771);
  nand GNAME4355(G4355,G21781,G1541);
  nand GNAME4356(G4356,G1543,G21590);
  nand GNAME4357(G4357,G1537,G8268);
  nand GNAME4358(G4358,G1538,G7477);
  nand GNAME4359(G4359,G1539,G7819);
  nand GNAME4360(G4360,G1540,G8785);
  nand GNAME4361(G4361,G21782,G1541);
  nand GNAME4362(G4362,G1543,G21591);
  nand GNAME4363(G4363,G1537,G8267);
  nand GNAME4364(G4364,G1538,G7476);
  nand GNAME4365(G4365,G1539,G7818);
  nand GNAME4366(G4366,G1540,G8704);
  nand GNAME4367(G4367,G21783,G1541);
  nand GNAME4368(G4368,G1543,G21592);
  nand GNAME4369(G4369,G1537,G8266);
  nand GNAME4370(G4370,G1538,G7475);
  nand GNAME4371(G4371,G1539,G7817);
  nand GNAME4372(G4372,G1540,G8705);
  nand GNAME4373(G4373,G21784,G1541);
  nand GNAME4374(G4374,G1543,G21593);
  nand GNAME4375(G4375,G1537,G8265);
  nand GNAME4376(G4376,G1538,G7474);
  nand GNAME4377(G4377,G1539,G7816);
  nand GNAME4378(G4378,G1540,G8761);
  nand GNAME4379(G4379,G21785,G1541);
  nand GNAME4380(G4380,G1543,G21594);
  nand GNAME4381(G4381,G1537,G8264);
  nand GNAME4382(G4382,G1538,G7473);
  nand GNAME4383(G4383,G1539,G7815);
  nand GNAME4384(G4384,G1540,G8706);
  nand GNAME4385(G4385,G21786,G1541);
  nand GNAME4386(G4386,G1543,G21595);
  nand GNAME4387(G4387,G1537,G8263);
  nand GNAME4388(G4388,G1538,G7472);
  nand GNAME4389(G4389,G1539,G7814);
  nand GNAME4390(G4390,G1540,G8707);
  nand GNAME4391(G4391,G21787,G1541);
  nand GNAME4392(G4392,G1543,G21596);
  nand GNAME4393(G4393,G1537,G8209);
  nand GNAME4394(G4394,G1538,G7441);
  nand GNAME4395(G4395,G1539,G7777);
  nand GNAME4396(G4396,G1540,G8760);
  nand GNAME4397(G4397,G21788,G1541);
  nand GNAME4398(G4398,G1543,G21597);
  nand GNAME4399(G4399,G1537,G8210);
  nand GNAME4400(G4400,G1538,G7442);
  nand GNAME4401(G4401,G1539,G7778);
  nand GNAME4402(G4402,G1540,G8770);
  nand GNAME4403(G4403,G21789,G1541);
  nand GNAME4404(G4404,G1543,G21598);
  nand GNAME4405(G4405,G2615,G1208,G1269);
  not GNAME4406(G4406,G1722);
  nand GNAME4407(G4407,G7809,G1546);
  nand GNAME4408(G4408,G21758,G1547);
  nand GNAME4409(G4409,G7467,G1548);
  nand GNAME4410(G4410,G8258,G1549);
  nand GNAME4411(G4411,G1550,G21599);
  nand GNAME4412(G4412,G7824,G1546);
  nand GNAME4413(G4413,G21759,G1547);
  nand GNAME4414(G4414,G7482,G1548);
  nand GNAME4415(G4415,G8273,G1549);
  nand GNAME4416(G4416,G1550,G21600);
  nand GNAME4417(G4417,G7776,G1546);
  nand GNAME4418(G4418,G21760,G1547);
  nand GNAME4419(G4419,G7440,G1548);
  nand GNAME4420(G4420,G8208,G1549);
  nand GNAME4421(G4421,G1550,G21601);
  nand GNAME4422(G4422,G7779,G1546);
  nand GNAME4423(G4423,G21761,G1547);
  nand GNAME4424(G4424,G7443,G1548);
  nand GNAME4425(G4425,G8211,G1549);
  nand GNAME4426(G4426,G1550,G21602);
  nand GNAME4427(G4427,G7813,G1546);
  nand GNAME4428(G4428,G21762,G1547);
  nand GNAME4429(G4429,G7471,G1548);
  nand GNAME4430(G4430,G8262,G1549);
  nand GNAME4431(G4431,G1550,G21603);
  nand GNAME4432(G4432,G7812,G1546);
  nand GNAME4433(G4433,G21763,G1547);
  nand GNAME4434(G4434,G7470,G1548);
  nand GNAME4435(G4435,G8261,G1549);
  nand GNAME4436(G4436,G1550,G21604);
  nand GNAME4437(G4437,G7780,G1546);
  nand GNAME4438(G4438,G21764,G1547);
  nand GNAME4439(G4439,G7444,G1548);
  nand GNAME4440(G4440,G8212,G1549);
  nand GNAME4441(G4441,G1550,G21605);
  nand GNAME4442(G4442,G7781,G1546);
  nand GNAME4443(G4443,G21765,G1547);
  nand GNAME4444(G4444,G7445,G1548);
  nand GNAME4445(G4445,G8213,G1549);
  nand GNAME4446(G4446,G1550,G21606);
  nand GNAME4447(G4447,G7811,G1546);
  nand GNAME4448(G4448,G21766,G1547);
  nand GNAME4449(G4449,G7469,G1548);
  nand GNAME4450(G4450,G8260,G1549);
  nand GNAME4451(G4451,G1550,G21607);
  nand GNAME4452(G4452,G7810,G1546);
  nand GNAME4453(G4453,G21767,G1547);
  nand GNAME4454(G4454,G7468,G1548);
  nand GNAME4455(G4455,G8259,G1549);
  nand GNAME4456(G4456,G1550,G21608);
  nand GNAME4457(G4457,G7773,G1546);
  nand GNAME4458(G4458,G21768,G1547);
  nand GNAME4459(G4459,G7437,G1548);
  nand GNAME4460(G4460,G8205,G1549);
  nand GNAME4461(G4461,G1550,G21609);
  nand GNAME4462(G4462,G7774,G1546);
  nand GNAME4463(G4463,G21769,G1547);
  nand GNAME4464(G4464,G7438,G1548);
  nand GNAME4465(G4465,G8206,G1549);
  nand GNAME4466(G4466,G1550,G21610);
  nand GNAME4467(G4467,G7831,G1546);
  nand GNAME4468(G4468,G21770,G1547);
  nand GNAME4469(G4469,G7489,G1548);
  nand GNAME4470(G4470,G8280,G1549);
  nand GNAME4471(G4471,G1550,G21611);
  nand GNAME4472(G4472,G7830,G1546);
  nand GNAME4473(G4473,G21771,G1547);
  nand GNAME4474(G4474,G7488,G1548);
  nand GNAME4475(G4475,G8279,G1549);
  nand GNAME4476(G4476,G1550,G21612);
  nand GNAME4477(G4477,G7775,G1546);
  nand GNAME4478(G4478,G21772,G1547);
  nand GNAME4479(G4479,G7439,G1548);
  nand GNAME4480(G4480,G8207,G1549);
  nand GNAME4481(G4481,G1550,G21613);
  nand GNAME4482(G4482,G7829,G1546);
  nand GNAME4483(G4483,G21773,G1547);
  nand GNAME4484(G4484,G7487,G1548);
  nand GNAME4485(G4485,G8278,G1549);
  nand GNAME4486(G4486,G1550,G21614);
  nand GNAME4487(G4487,G7828,G1546);
  nand GNAME4488(G4488,G21774,G1547);
  nand GNAME4489(G4489,G7486,G1548);
  nand GNAME4490(G4490,G8277,G1549);
  nand GNAME4491(G4491,G1550,G21615);
  nand GNAME4492(G4492,G7827,G1546);
  nand GNAME4493(G4493,G21775,G1547);
  nand GNAME4494(G4494,G7485,G1548);
  nand GNAME4495(G4495,G8276,G1549);
  nand GNAME4496(G4496,G1550,G21616);
  nand GNAME4497(G4497,G7826,G1546);
  nand GNAME4498(G4498,G21776,G1547);
  nand GNAME4499(G4499,G7484,G1548);
  nand GNAME4500(G4500,G8275,G1549);
  nand GNAME4501(G4501,G1550,G21617);
  nand GNAME4502(G4502,G7825,G1546);
  nand GNAME4503(G4503,G21777,G1547);
  nand GNAME4504(G4504,G7483,G1548);
  nand GNAME4505(G4505,G8274,G1549);
  nand GNAME4506(G4506,G1550,G21618);
  nand GNAME4507(G4507,G7823,G1546);
  nand GNAME4508(G4508,G21778,G1547);
  nand GNAME4509(G4509,G7481,G1548);
  nand GNAME4510(G4510,G8272,G1549);
  nand GNAME4511(G4511,G1550,G21619);
  nand GNAME4512(G4512,G7822,G1546);
  nand GNAME4513(G4513,G21779,G1547);
  nand GNAME4514(G4514,G7480,G1548);
  nand GNAME4515(G4515,G8271,G1549);
  nand GNAME4516(G4516,G1550,G21620);
  nand GNAME4517(G4517,G7821,G1546);
  nand GNAME4518(G4518,G21780,G1547);
  nand GNAME4519(G4519,G7479,G1548);
  nand GNAME4520(G4520,G8270,G1549);
  nand GNAME4521(G4521,G1550,G21621);
  nand GNAME4522(G4522,G7820,G1546);
  nand GNAME4523(G4523,G21781,G1547);
  nand GNAME4524(G4524,G7478,G1548);
  nand GNAME4525(G4525,G8269,G1549);
  nand GNAME4526(G4526,G1550,G21622);
  nand GNAME4527(G4527,G7819,G1546);
  nand GNAME4528(G4528,G21782,G1547);
  nand GNAME4529(G4529,G7477,G1548);
  nand GNAME4530(G4530,G8268,G1549);
  nand GNAME4531(G4531,G1550,G21623);
  nand GNAME4532(G4532,G7818,G1546);
  nand GNAME4533(G4533,G21783,G1547);
  nand GNAME4534(G4534,G7476,G1548);
  nand GNAME4535(G4535,G8267,G1549);
  nand GNAME4536(G4536,G1550,G21624);
  nand GNAME4537(G4537,G7817,G1546);
  nand GNAME4538(G4538,G21784,G1547);
  nand GNAME4539(G4539,G7475,G1548);
  nand GNAME4540(G4540,G8266,G1549);
  nand GNAME4541(G4541,G1550,G21625);
  nand GNAME4542(G4542,G7816,G1546);
  nand GNAME4543(G4543,G21785,G1547);
  nand GNAME4544(G4544,G7474,G1548);
  nand GNAME4545(G4545,G8265,G1549);
  nand GNAME4546(G4546,G1550,G21626);
  nand GNAME4547(G4547,G7815,G1546);
  nand GNAME4548(G4548,G21786,G1547);
  nand GNAME4549(G4549,G7473,G1548);
  nand GNAME4550(G4550,G8264,G1549);
  nand GNAME4551(G4551,G1550,G21627);
  nand GNAME4552(G4552,G7814,G1546);
  nand GNAME4553(G4553,G21787,G1547);
  nand GNAME4554(G4554,G7472,G1548);
  nand GNAME4555(G4555,G8263,G1549);
  nand GNAME4556(G4556,G1550,G21628);
  nand GNAME4557(G4557,G7777,G1546);
  nand GNAME4558(G4558,G21788,G1547);
  nand GNAME4559(G4559,G7441,G1548);
  nand GNAME4560(G4560,G8209,G1549);
  nand GNAME4561(G4561,G1550,G21629);
  nand GNAME4562(G4562,G7778,G1546);
  nand GNAME4563(G4563,G21789,G1547);
  nand GNAME4564(G4564,G7442,G1548);
  nand GNAME4565(G4565,G8210,G1549);
  nand GNAME4566(G4566,G1550,G21630);
  nand GNAME4567(G4567,G1506,G2320,G7326);
  or GNAME4568(G4568,G2332,G1552);
  nand GNAME4569(G4569,G1553,G21709);
  nand GNAME4570(G4570,G1554,G17);
  nand GNAME4571(G4571,G1555,G21631);
  nand GNAME4572(G4572,G1553,G21708);
  nand GNAME4573(G4573,G1555,G21632);
  nand GNAME4574(G4574,G1553,G21707);
  nand GNAME4575(G4575,G1555,G21633);
  nand GNAME4576(G4576,G1553,G21706);
  nand GNAME4577(G4577,G1555,G21634);
  nand GNAME4578(G4578,G1553,G21705);
  nand GNAME4579(G4579,G1555,G21635);
  nand GNAME4580(G4580,G1553,G21704);
  nand GNAME4581(G4581,G1555,G21636);
  nand GNAME4582(G4582,G1553,G21703);
  nand GNAME4583(G4583,G1555,G21637);
  nand GNAME4584(G4584,G1553,G21702);
  nand GNAME4585(G4585,G1555,G21638);
  nand GNAME4586(G4586,G1553,G21701);
  nand GNAME4587(G4587,G1555,G21639);
  nand GNAME4588(G4588,G1553,G21700);
  nand GNAME4589(G4589,G1555,G21640);
  nand GNAME4590(G4590,G1553,G21699);
  nand GNAME4591(G4591,G1555,G21641);
  nand GNAME4592(G4592,G1553,G21698);
  nand GNAME4593(G4593,G1555,G21642);
  nand GNAME4594(G4594,G1553,G21697);
  nand GNAME4595(G4595,G1555,G21643);
  nand GNAME4596(G4596,G1553,G21696);
  nand GNAME4597(G4597,G1555,G21644);
  nand GNAME4598(G4598,G1553,G21695);
  nand GNAME4599(G4599,G1555,G21645);
  nand GNAME4600(G4600,G1553,G21694);
  nand GNAME4601(G4601,G1555,G21646);
  nand GNAME4602(G4602,G1553,G21724);
  nand GNAME4603(G4603,G1554,G18);
  nand GNAME4604(G4604,G1555,G21647);
  nand GNAME4605(G4605,G1553,G21723);
  nand GNAME4606(G4606,G1554,G19);
  nand GNAME4607(G4607,G1555,G21648);
  nand GNAME4608(G4608,G1553,G21722);
  nand GNAME4609(G4609,G1554,G20);
  nand GNAME4610(G4610,G1555,G21649);
  nand GNAME4611(G4611,G1553,G21721);
  nand GNAME4612(G4612,G1554,G21);
  nand GNAME4613(G4613,G1555,G21650);
  nand GNAME4614(G4614,G1553,G21720);
  nand GNAME4615(G4615,G1554,G22);
  nand GNAME4616(G4616,G1555,G21651);
  nand GNAME4617(G4617,G1553,G21719);
  nand GNAME4618(G4618,G1554,G23);
  nand GNAME4619(G4619,G1555,G21652);
  nand GNAME4620(G4620,G1553,G21718);
  nand GNAME4621(G4621,G1554,G24);
  nand GNAME4622(G4622,G1555,G21653);
  nand GNAME4623(G4623,G1553,G21717);
  nand GNAME4624(G4624,G25,G1554);
  nand GNAME4625(G4625,G1555,G21654);
  nand GNAME4626(G4626,G1553,G21716);
  nand GNAME4627(G4627,G26,G1554);
  nand GNAME4628(G4628,G1555,G21655);
  nand GNAME4629(G4629,G1553,G21715);
  nand GNAME4630(G4630,G27,G1554);
  nand GNAME4631(G4631,G1555,G21656);
  nand GNAME4632(G4632,G1553,G21714);
  nand GNAME4633(G4633,G28,G1554);
  nand GNAME4634(G4634,G1555,G21657);
  nand GNAME4635(G4635,G1553,G21713);
  nand GNAME4636(G4636,G29,G1554);
  nand GNAME4637(G4637,G1555,G21658);
  nand GNAME4638(G4638,G1553,G21712);
  nand GNAME4639(G4639,G30,G1554);
  nand GNAME4640(G4640,G1555,G21659);
  nand GNAME4641(G4641,G1553,G21711);
  nand GNAME4642(G4642,G31,G1554);
  nand GNAME4643(G4643,G1555,G21660);
  nand GNAME4644(G4644,G1553,G21710);
  nand GNAME4645(G4645,G32,G1554);
  nand GNAME4646(G4646,G1555,G21661);
  nand GNAME4647(G4647,G2460,G2308);
  or GNAME4648(G4648,G21392,G1558);
  nand GNAME4649(G4649,G4647,G4648);
  nand GNAME4650(G4650,G1283,G4649,G7326);
  nand GNAME4651(G4651,G21427,G1292);
  nand GNAME4652(G4652,G21646,G1559);
  nand GNAME4653(G4653,G21694,G1560);
  nand GNAME4654(G4654,G1561,G21662);
  nand GNAME4655(G4655,G21645,G1559);
  nand GNAME4656(G4656,G21695,G1560);
  nand GNAME4657(G4657,G1561,G21663);
  nand GNAME4658(G4658,G21644,G1559);
  nand GNAME4659(G4659,G21696,G1560);
  nand GNAME4660(G4660,G1561,G21664);
  nand GNAME4661(G4661,G21643,G1559);
  nand GNAME4662(G4662,G21697,G1560);
  nand GNAME4663(G4663,G1561,G21665);
  nand GNAME4664(G4664,G21642,G1559);
  nand GNAME4665(G4665,G21698,G1560);
  nand GNAME4666(G4666,G1561,G21666);
  nand GNAME4667(G4667,G21641,G1559);
  nand GNAME4668(G4668,G21699,G1560);
  nand GNAME4669(G4669,G1561,G21667);
  nand GNAME4670(G4670,G21640,G1559);
  nand GNAME4671(G4671,G21700,G1560);
  nand GNAME4672(G4672,G1561,G21668);
  nand GNAME4673(G4673,G21639,G1559);
  nand GNAME4674(G4674,G21701,G1560);
  nand GNAME4675(G4675,G1561,G21669);
  nand GNAME4676(G4676,G21638,G1559);
  nand GNAME4677(G4677,G21702,G1560);
  nand GNAME4678(G4678,G1561,G21670);
  nand GNAME4679(G4679,G21637,G1559);
  nand GNAME4680(G4680,G21703,G1560);
  nand GNAME4681(G4681,G1561,G21671);
  nand GNAME4682(G4682,G21636,G1559);
  nand GNAME4683(G4683,G21704,G1560);
  nand GNAME4684(G4684,G1561,G21672);
  nand GNAME4685(G4685,G21635,G1559);
  nand GNAME4686(G4686,G21705,G1560);
  nand GNAME4687(G4687,G1561,G21673);
  nand GNAME4688(G4688,G21634,G1559);
  nand GNAME4689(G4689,G21706,G1560);
  nand GNAME4690(G4690,G1561,G21674);
  nand GNAME4691(G4691,G21633,G1559);
  nand GNAME4692(G4692,G21707,G1560);
  nand GNAME4693(G4693,G1561,G21675);
  nand GNAME4694(G4694,G21632,G1559);
  nand GNAME4695(G4695,G21708,G1560);
  nand GNAME4696(G4696,G1561,G21676);
  nand GNAME4697(G4697,G21631,G1559);
  nand GNAME4698(G4698,G21709,G1560);
  nand GNAME4699(G4699,G1561,G21677);
  nand GNAME4700(G4700,G21710,G1562);
  nand GNAME4701(G4701,G21661,G1559);
  nand GNAME4702(G4702,G1561,G21678);
  nand GNAME4703(G4703,G21711,G1562);
  nand GNAME4704(G4704,G21660,G1559);
  nand GNAME4705(G4705,G1561,G21679);
  nand GNAME4706(G4706,G21712,G1562);
  nand GNAME4707(G4707,G21659,G1559);
  nand GNAME4708(G4708,G1561,G21680);
  nand GNAME4709(G4709,G21713,G1562);
  nand GNAME4710(G4710,G21658,G1559);
  nand GNAME4711(G4711,G1561,G21681);
  nand GNAME4712(G4712,G21714,G1562);
  nand GNAME4713(G4713,G21657,G1559);
  nand GNAME4714(G4714,G1561,G21682);
  nand GNAME4715(G4715,G21715,G1562);
  nand GNAME4716(G4716,G21656,G1559);
  nand GNAME4717(G4717,G1561,G21683);
  nand GNAME4718(G4718,G21716,G1562);
  nand GNAME4719(G4719,G21655,G1559);
  nand GNAME4720(G4720,G1561,G21684);
  nand GNAME4721(G4721,G21717,G1562);
  nand GNAME4722(G4722,G21654,G1559);
  nand GNAME4723(G4723,G1561,G21685);
  nand GNAME4724(G4724,G21718,G1562);
  nand GNAME4725(G4725,G21653,G1559);
  nand GNAME4726(G4726,G1561,G21686);
  nand GNAME4727(G4727,G21719,G1562);
  nand GNAME4728(G4728,G21652,G1559);
  nand GNAME4729(G4729,G1561,G21687);
  nand GNAME4730(G4730,G21720,G1562);
  nand GNAME4731(G4731,G21651,G1559);
  nand GNAME4732(G4732,G1561,G21688);
  nand GNAME4733(G4733,G21721,G1562);
  nand GNAME4734(G4734,G21650,G1559);
  nand GNAME4735(G4735,G1561,G21689);
  nand GNAME4736(G4736,G21722,G1562);
  nand GNAME4737(G4737,G21649,G1559);
  nand GNAME4738(G4738,G1561,G21690);
  nand GNAME4739(G4739,G21723,G1562);
  nand GNAME4740(G4740,G21648,G1559);
  nand GNAME4741(G4741,G1561,G21691);
  nand GNAME4742(G4742,G21724,G1562);
  nand GNAME4743(G4743,G21647,G1559);
  nand GNAME4744(G4744,G1561,G21692);
  nand GNAME4745(G4745,G1202,G1564);
  nand GNAME4746(G4746,G4745,G1713);
  nand GNAME4747(G4747,G4746,G7326);
  nand GNAME4748(G4748,G4747,G1723,G1552);
  nand GNAME4749(G4749,G32,G1566);
  nand GNAME4750(G4750,G8258,G1567);
  nand GNAME4751(G4751,G7467,G1568);
  nand GNAME4752(G4752,G1565,G21694);
  nand GNAME4753(G4753,G31,G1566);
  nand GNAME4754(G4754,G8273,G1567);
  nand GNAME4755(G4755,G7482,G1568);
  nand GNAME4756(G4756,G1565,G21695);
  nand GNAME4757(G4757,G30,G1566);
  nand GNAME4758(G4758,G8208,G1567);
  nand GNAME4759(G4759,G7440,G1568);
  nand GNAME4760(G4760,G1565,G21696);
  nand GNAME4761(G4761,G29,G1566);
  nand GNAME4762(G4762,G8211,G1567);
  nand GNAME4763(G4763,G7443,G1568);
  nand GNAME4764(G4764,G1565,G21697);
  nand GNAME4765(G4765,G28,G1566);
  nand GNAME4766(G4766,G8262,G1567);
  nand GNAME4767(G4767,G7471,G1568);
  nand GNAME4768(G4768,G1565,G21698);
  nand GNAME4769(G4769,G27,G1566);
  nand GNAME4770(G4770,G8261,G1567);
  nand GNAME4771(G4771,G7470,G1568);
  nand GNAME4772(G4772,G1565,G21699);
  nand GNAME4773(G4773,G26,G1566);
  nand GNAME4774(G4774,G8212,G1567);
  nand GNAME4775(G4775,G7444,G1568);
  nand GNAME4776(G4776,G1565,G21700);
  nand GNAME4777(G4777,G25,G1566);
  nand GNAME4778(G4778,G8213,G1567);
  nand GNAME4779(G4779,G7445,G1568);
  nand GNAME4780(G4780,G1565,G21701);
  nand GNAME4781(G4781,G24,G1566);
  nand GNAME4782(G4782,G8260,G1567);
  nand GNAME4783(G4783,G7469,G1568);
  nand GNAME4784(G4784,G1565,G21702);
  nand GNAME4785(G4785,G23,G1566);
  nand GNAME4786(G4786,G8259,G1567);
  nand GNAME4787(G4787,G7468,G1568);
  nand GNAME4788(G4788,G1565,G21703);
  nand GNAME4789(G4789,G22,G1566);
  nand GNAME4790(G4790,G8205,G1567);
  nand GNAME4791(G4791,G7437,G1568);
  nand GNAME4792(G4792,G1565,G21704);
  nand GNAME4793(G4793,G21,G1566);
  nand GNAME4794(G4794,G8206,G1567);
  nand GNAME4795(G4795,G7438,G1568);
  nand GNAME4796(G4796,G1565,G21705);
  nand GNAME4797(G4797,G20,G1566);
  nand GNAME4798(G4798,G8280,G1567);
  nand GNAME4799(G4799,G7489,G1568);
  nand GNAME4800(G4800,G1565,G21706);
  nand GNAME4801(G4801,G19,G1566);
  nand GNAME4802(G4802,G8279,G1567);
  nand GNAME4803(G4803,G7488,G1568);
  nand GNAME4804(G4804,G1565,G21707);
  nand GNAME4805(G4805,G18,G1566);
  nand GNAME4806(G4806,G8207,G1567);
  nand GNAME4807(G4807,G7439,G1568);
  nand GNAME4808(G4808,G1565,G21708);
  nand GNAME4809(G4809,G17,G1566);
  nand GNAME4810(G4810,G8278,G1567);
  nand GNAME4811(G4811,G7487,G1568);
  nand GNAME4812(G4812,G1565,G21709);
  nand GNAME4813(G4813,G32,G1569);
  nand GNAME4814(G4814,G16,G1570);
  nand GNAME4815(G4815,G8277,G1567);
  nand GNAME4816(G4816,G7486,G1568);
  nand GNAME4817(G4817,G1565,G21710);
  nand GNAME4818(G4818,G31,G1569);
  nand GNAME4819(G4819,G15,G1570);
  nand GNAME4820(G4820,G8276,G1567);
  nand GNAME4821(G4821,G7485,G1568);
  nand GNAME4822(G4822,G1565,G21711);
  nand GNAME4823(G4823,G30,G1569);
  nand GNAME4824(G4824,G14,G1570);
  nand GNAME4825(G4825,G8275,G1567);
  nand GNAME4826(G4826,G7484,G1568);
  nand GNAME4827(G4827,G1565,G21712);
  nand GNAME4828(G4828,G29,G1569);
  nand GNAME4829(G4829,G13,G1570);
  nand GNAME4830(G4830,G8274,G1567);
  nand GNAME4831(G4831,G7483,G1568);
  nand GNAME4832(G4832,G1565,G21713);
  nand GNAME4833(G4833,G28,G1569);
  nand GNAME4834(G4834,G12,G1570);
  nand GNAME4835(G4835,G8272,G1567);
  nand GNAME4836(G4836,G7481,G1568);
  nand GNAME4837(G4837,G1565,G21714);
  nand GNAME4838(G4838,G27,G1569);
  nand GNAME4839(G4839,G11,G1570);
  nand GNAME4840(G4840,G8271,G1567);
  nand GNAME4841(G4841,G7480,G1568);
  nand GNAME4842(G4842,G1565,G21715);
  nand GNAME4843(G4843,G26,G1569);
  nand GNAME4844(G4844,G10,G1570);
  nand GNAME4845(G4845,G8270,G1567);
  nand GNAME4846(G4846,G7479,G1568);
  nand GNAME4847(G4847,G1565,G21716);
  nand GNAME4848(G4848,G25,G1569);
  nand GNAME4849(G4849,G9,G1570);
  nand GNAME4850(G4850,G8269,G1567);
  nand GNAME4851(G4851,G7478,G1568);
  nand GNAME4852(G4852,G1565,G21717);
  nand GNAME4853(G4853,G24,G1569);
  nand GNAME4854(G4854,G8,G1570);
  nand GNAME4855(G4855,G8268,G1567);
  nand GNAME4856(G4856,G7477,G1568);
  nand GNAME4857(G4857,G1565,G21718);
  nand GNAME4858(G4858,G23,G1569);
  nand GNAME4859(G4859,G7,G1570);
  nand GNAME4860(G4860,G8267,G1567);
  nand GNAME4861(G4861,G7476,G1568);
  nand GNAME4862(G4862,G1565,G21719);
  nand GNAME4863(G4863,G22,G1569);
  nand GNAME4864(G4864,G6,G1570);
  nand GNAME4865(G4865,G8266,G1567);
  nand GNAME4866(G4866,G7475,G1568);
  nand GNAME4867(G4867,G1565,G21720);
  nand GNAME4868(G4868,G21,G1569);
  nand GNAME4869(G4869,G5,G1570);
  nand GNAME4870(G4870,G8265,G1567);
  nand GNAME4871(G4871,G7474,G1568);
  nand GNAME4872(G4872,G1565,G21721);
  nand GNAME4873(G4873,G20,G1569);
  nand GNAME4874(G4874,G4,G1570);
  nand GNAME4875(G4875,G8264,G1567);
  nand GNAME4876(G4876,G7473,G1568);
  nand GNAME4877(G4877,G1565,G21722);
  nand GNAME4878(G4878,G19,G1569);
  nand GNAME4879(G4879,G3,G1570);
  nand GNAME4880(G4880,G8263,G1567);
  nand GNAME4881(G4881,G7472,G1568);
  nand GNAME4882(G4882,G1565,G21723);
  nand GNAME4883(G4883,G18,G1569);
  nand GNAME4884(G4884,G2,G1570);
  nand GNAME4885(G4885,G8209,G1567);
  nand GNAME4886(G4886,G7441,G1568);
  nand GNAME4887(G4887,G1565,G21724);
  nand GNAME4888(G4888,G1,G1570);
  nand GNAME4889(G4889,G7442,G1568);
  nand GNAME4890(G4890,G1565,G21725);
  nand GNAME4891(G4891,G7326,G1571);
  nand GNAME4892(G4892,G4891,G2299);
  nand GNAME4893(G4893,G7809,G1574);
  nand GNAME4894(G4894,G7467,G1575);
  nand GNAME4895(G4895,G1573,G21726);
  nand GNAME4896(G4896,G7824,G1574);
  nand GNAME4897(G4897,G7482,G1575);
  nand GNAME4898(G4898,G1573,G21727);
  nand GNAME4899(G4899,G7776,G1574);
  nand GNAME4900(G4900,G7440,G1575);
  nand GNAME4901(G4901,G1573,G21728);
  nand GNAME4902(G4902,G7779,G1574);
  nand GNAME4903(G4903,G7443,G1575);
  nand GNAME4904(G4904,G1573,G21729);
  nand GNAME4905(G4905,G7813,G1574);
  nand GNAME4906(G4906,G7471,G1575);
  nand GNAME4907(G4907,G1573,G21730);
  nand GNAME4908(G4908,G7812,G1574);
  nand GNAME4909(G4909,G7470,G1575);
  nand GNAME4910(G4910,G1573,G21731);
  nand GNAME4911(G4911,G7780,G1574);
  nand GNAME4912(G4912,G7444,G1575);
  nand GNAME4913(G4913,G1573,G21732);
  nand GNAME4914(G4914,G7781,G1574);
  nand GNAME4915(G4915,G7445,G1575);
  nand GNAME4916(G4916,G1573,G21733);
  nand GNAME4917(G4917,G7811,G1574);
  nand GNAME4918(G4918,G7469,G1575);
  nand GNAME4919(G4919,G1573,G21734);
  nand GNAME4920(G4920,G7810,G1574);
  nand GNAME4921(G4921,G7468,G1575);
  nand GNAME4922(G4922,G1573,G21735);
  nand GNAME4923(G4923,G7773,G1574);
  nand GNAME4924(G4924,G7437,G1575);
  nand GNAME4925(G4925,G1573,G21736);
  nand GNAME4926(G4926,G7774,G1574);
  nand GNAME4927(G4927,G7438,G1575);
  nand GNAME4928(G4928,G1573,G21737);
  nand GNAME4929(G4929,G7831,G1574);
  nand GNAME4930(G4930,G7489,G1575);
  nand GNAME4931(G4931,G1573,G21738);
  nand GNAME4932(G4932,G7830,G1574);
  nand GNAME4933(G4933,G7488,G1575);
  nand GNAME4934(G4934,G1573,G21739);
  nand GNAME4935(G4935,G7775,G1574);
  nand GNAME4936(G4936,G7439,G1575);
  nand GNAME4937(G4937,G1573,G21740);
  nand GNAME4938(G4938,G7829,G1574);
  nand GNAME4939(G4939,G7487,G1575);
  nand GNAME4940(G4940,G1573,G21741);
  nand GNAME4941(G4941,G7828,G1574);
  nand GNAME4942(G4942,G7486,G1575);
  nand GNAME4943(G4943,G1573,G21742);
  nand GNAME4944(G4944,G7827,G1574);
  nand GNAME4945(G4945,G7485,G1575);
  nand GNAME4946(G4946,G1573,G21743);
  nand GNAME4947(G4947,G7826,G1574);
  nand GNAME4948(G4948,G7484,G1575);
  nand GNAME4949(G4949,G1573,G21744);
  nand GNAME4950(G4950,G7825,G1574);
  nand GNAME4951(G4951,G7483,G1575);
  nand GNAME4952(G4952,G1573,G21745);
  nand GNAME4953(G4953,G7823,G1574);
  nand GNAME4954(G4954,G7481,G1575);
  nand GNAME4955(G4955,G1573,G21746);
  nand GNAME4956(G4956,G7822,G1574);
  nand GNAME4957(G4957,G7480,G1575);
  nand GNAME4958(G4958,G1573,G21747);
  nand GNAME4959(G4959,G7821,G1574);
  nand GNAME4960(G4960,G7479,G1575);
  nand GNAME4961(G4961,G1573,G21748);
  nand GNAME4962(G4962,G7820,G1574);
  nand GNAME4963(G4963,G7478,G1575);
  nand GNAME4964(G4964,G1573,G21749);
  nand GNAME4965(G4965,G7819,G1574);
  nand GNAME4966(G4966,G7477,G1575);
  nand GNAME4967(G4967,G1573,G21750);
  nand GNAME4968(G4968,G7818,G1574);
  nand GNAME4969(G4969,G7476,G1575);
  nand GNAME4970(G4970,G1573,G21751);
  nand GNAME4971(G4971,G7817,G1574);
  nand GNAME4972(G4972,G7475,G1575);
  nand GNAME4973(G4973,G1573,G21752);
  nand GNAME4974(G4974,G7816,G1574);
  nand GNAME4975(G4975,G7474,G1575);
  nand GNAME4976(G4976,G1573,G21753);
  nand GNAME4977(G4977,G7815,G1574);
  nand GNAME4978(G4978,G7473,G1575);
  nand GNAME4979(G4979,G1573,G21754);
  nand GNAME4980(G4980,G7814,G1574);
  nand GNAME4981(G4981,G7472,G1575);
  nand GNAME4982(G4982,G1573,G21755);
  nand GNAME4983(G4983,G7777,G1574);
  nand GNAME4984(G4984,G7441,G1575);
  nand GNAME4985(G4985,G1573,G21756);
  nand GNAME4986(G4986,G7442,G1575);
  nand GNAME4987(G4987,G1573,G21757);
  nand GNAME4988(G4988,G1251,G1299,G2511,G1240,G21426);
  nand GNAME4989(G4989,G2320,G1506);
  nand GNAME4990(G4990,G2297,G1283,G8101);
  or GNAME4991(G4991,G1588,G1282);
  not GNAME4992(G4992,G1583);
  or GNAME4993(G4993,G2329,G1209,G1245);
  nand GNAME4994(G4994,G21427,G7442);
  nand GNAME4995(G4995,G21426,G1511);
  nand GNAME4996(G4996,G4995,G1580);
  or GNAME4997(G4997,G35,G21797);
  nand GNAME4998(G4998,G6742,G8258);
  nand GNAME4999(G4999,G6741,G7467);
  nand GNAME5000(G5000,G6740,G21726);
  nand GNAME5001(G5001,G7809,G1581);
  nand GNAME5002(G5002,G21599,G1582);
  nand GNAME5003(G5003,G21758,G4992);
  nand GNAME5004(G5004,G6742,G8273);
  nand GNAME5005(G5005,G6741,G7482);
  nand GNAME5006(G5006,G6740,G21727);
  nand GNAME5007(G5007,G7824,G1581);
  nand GNAME5008(G5008,G21600,G1582);
  nand GNAME5009(G5009,G21759,G4992);
  nand GNAME5010(G5010,G6742,G8208);
  nand GNAME5011(G5011,G6741,G7440);
  nand GNAME5012(G5012,G6740,G21728);
  nand GNAME5013(G5013,G7776,G1581);
  nand GNAME5014(G5014,G21601,G1582);
  nand GNAME5015(G5015,G21760,G4992);
  nand GNAME5016(G5016,G6742,G8211);
  nand GNAME5017(G5017,G6741,G7443);
  nand GNAME5018(G5018,G6740,G21729);
  nand GNAME5019(G5019,G7779,G1581);
  nand GNAME5020(G5020,G21602,G1582);
  nand GNAME5021(G5021,G21761,G4992);
  nand GNAME5022(G5022,G6742,G8262);
  nand GNAME5023(G5023,G6741,G7471);
  nand GNAME5024(G5024,G6740,G21730);
  nand GNAME5025(G5025,G7813,G1581);
  nand GNAME5026(G5026,G21603,G1582);
  nand GNAME5027(G5027,G21762,G4992);
  nand GNAME5028(G5028,G6742,G8261);
  nand GNAME5029(G5029,G6741,G7470);
  nand GNAME5030(G5030,G6740,G21731);
  nand GNAME5031(G5031,G7812,G1581);
  nand GNAME5032(G5032,G21604,G1582);
  nand GNAME5033(G5033,G21763,G4992);
  nand GNAME5034(G5034,G8212,G1584);
  nand GNAME5035(G5035,G6741,G7444);
  nand GNAME5036(G5036,G6740,G21732);
  nand GNAME5037(G5037,G7780,G1585);
  nand GNAME5038(G5038,G21605,G1582);
  nand GNAME5039(G5039,G21764,G4992);
  nand GNAME5040(G5040,G8213,G1584);
  nand GNAME5041(G5041,G6741,G7445);
  nand GNAME5042(G5042,G6740,G21733);
  nand GNAME5043(G5043,G7781,G1585);
  nand GNAME5044(G5044,G21606,G1582);
  nand GNAME5045(G5045,G21765,G4992);
  nand GNAME5046(G5046,G8260,G1584);
  nand GNAME5047(G5047,G6741,G7469);
  nand GNAME5048(G5048,G6740,G21734);
  nand GNAME5049(G5049,G7811,G1585);
  nand GNAME5050(G5050,G21607,G1582);
  nand GNAME5051(G5051,G21766,G4992);
  nand GNAME5052(G5052,G8259,G1584);
  nand GNAME5053(G5053,G6741,G7468);
  nand GNAME5054(G5054,G6740,G21735);
  nand GNAME5055(G5055,G7810,G1585);
  nand GNAME5056(G5056,G21608,G1582);
  nand GNAME5057(G5057,G21767,G4992);
  nand GNAME5058(G5058,G8205,G1584);
  nand GNAME5059(G5059,G6741,G7437);
  nand GNAME5060(G5060,G6740,G21736);
  nand GNAME5061(G5061,G7773,G1585);
  nand GNAME5062(G5062,G21609,G1582);
  nand GNAME5063(G5063,G21768,G4992);
  nand GNAME5064(G5064,G8206,G1584);
  nand GNAME5065(G5065,G6741,G7438);
  nand GNAME5066(G5066,G6740,G21737);
  nand GNAME5067(G5067,G7774,G1585);
  nand GNAME5068(G5068,G21610,G1582);
  nand GNAME5069(G5069,G21769,G4992);
  nand GNAME5070(G5070,G8280,G1584);
  nand GNAME5071(G5071,G6741,G7489);
  nand GNAME5072(G5072,G6740,G21738);
  nand GNAME5073(G5073,G7831,G1585);
  nand GNAME5074(G5074,G21611,G1582);
  nand GNAME5075(G5075,G21770,G4992);
  nand GNAME5076(G5076,G8279,G1584);
  nand GNAME5077(G5077,G6741,G7488);
  nand GNAME5078(G5078,G6740,G21739);
  nand GNAME5079(G5079,G7830,G1585);
  nand GNAME5080(G5080,G21612,G1582);
  nand GNAME5081(G5081,G21771,G4992);
  nand GNAME5082(G5082,G8207,G1584);
  nand GNAME5083(G5083,G6741,G7439);
  nand GNAME5084(G5084,G6740,G21740);
  nand GNAME5085(G5085,G7775,G1585);
  nand GNAME5086(G5086,G21613,G1582);
  nand GNAME5087(G5087,G21772,G4992);
  nand GNAME5088(G5088,G8278,G1584);
  nand GNAME5089(G5089,G6741,G7487);
  nand GNAME5090(G5090,G6740,G21741);
  nand GNAME5091(G5091,G7829,G1585);
  nand GNAME5092(G5092,G21614,G1582);
  nand GNAME5093(G5093,G21773,G4992);
  nand GNAME5094(G5094,G8277,G1584);
  nand GNAME5095(G5095,G6741,G7486);
  nand GNAME5096(G5096,G6740,G21742);
  nand GNAME5097(G5097,G7828,G1585);
  nand GNAME5098(G5098,G21615,G1582);
  nand GNAME5099(G5099,G21774,G4992);
  nand GNAME5100(G5100,G8276,G1584);
  nand GNAME5101(G5101,G6741,G7485);
  nand GNAME5102(G5102,G6740,G21743);
  nand GNAME5103(G5103,G7827,G1585);
  nand GNAME5104(G5104,G21616,G1582);
  nand GNAME5105(G5105,G21775,G4992);
  nand GNAME5106(G5106,G8275,G1584);
  nand GNAME5107(G5107,G6741,G7484);
  nand GNAME5108(G5108,G6740,G21744);
  nand GNAME5109(G5109,G7826,G1585);
  nand GNAME5110(G5110,G21617,G1582);
  nand GNAME5111(G5111,G21776,G4992);
  nand GNAME5112(G5112,G8274,G1584);
  nand GNAME5113(G5113,G6741,G7483);
  nand GNAME5114(G5114,G6740,G21745);
  nand GNAME5115(G5115,G7825,G1585);
  nand GNAME5116(G5116,G21618,G1582);
  nand GNAME5117(G5117,G21777,G4992);
  nand GNAME5118(G5118,G8272,G1584);
  nand GNAME5119(G5119,G6741,G7481);
  nand GNAME5120(G5120,G6740,G21746);
  nand GNAME5121(G5121,G7823,G1585);
  nand GNAME5122(G5122,G21619,G1582);
  nand GNAME5123(G5123,G21778,G4992);
  nand GNAME5124(G5124,G8271,G1584);
  nand GNAME5125(G5125,G6741,G7480);
  nand GNAME5126(G5126,G6740,G21747);
  nand GNAME5127(G5127,G7822,G1585);
  nand GNAME5128(G5128,G21620,G1582);
  nand GNAME5129(G5129,G21779,G4992);
  nand GNAME5130(G5130,G8270,G1584);
  nand GNAME5131(G5131,G6741,G7479);
  nand GNAME5132(G5132,G6740,G21748);
  nand GNAME5133(G5133,G7821,G1585);
  nand GNAME5134(G5134,G21621,G1582);
  nand GNAME5135(G5135,G21780,G4992);
  nand GNAME5136(G5136,G8269,G1584);
  nand GNAME5137(G5137,G6741,G7478);
  nand GNAME5138(G5138,G6740,G21749);
  nand GNAME5139(G5139,G7820,G1585);
  nand GNAME5140(G5140,G21622,G1582);
  nand GNAME5141(G5141,G21781,G4992);
  nand GNAME5142(G5142,G8268,G1584);
  nand GNAME5143(G5143,G6741,G7477);
  nand GNAME5144(G5144,G6740,G21750);
  nand GNAME5145(G5145,G7819,G1585);
  nand GNAME5146(G5146,G21623,G1582);
  nand GNAME5147(G5147,G21782,G4992);
  nand GNAME5148(G5148,G8267,G1584);
  nand GNAME5149(G5149,G6741,G7476);
  nand GNAME5150(G5150,G6740,G21751);
  nand GNAME5151(G5151,G7818,G1585);
  nand GNAME5152(G5152,G21624,G1582);
  nand GNAME5153(G5153,G21783,G4992);
  nand GNAME5154(G5154,G8266,G1584);
  nand GNAME5155(G5155,G6741,G7475);
  nand GNAME5156(G5156,G6740,G21752);
  nand GNAME5157(G5157,G7817,G1585);
  nand GNAME5158(G5158,G21625,G1582);
  nand GNAME5159(G5159,G21784,G4992);
  nand GNAME5160(G5160,G8265,G1584);
  nand GNAME5161(G5161,G6741,G7474);
  nand GNAME5162(G5162,G6740,G21753);
  nand GNAME5163(G5163,G7816,G1585);
  nand GNAME5164(G5164,G21626,G1582);
  nand GNAME5165(G5165,G21785,G4992);
  nand GNAME5166(G5166,G8264,G1584);
  nand GNAME5167(G5167,G6741,G7473);
  nand GNAME5168(G5168,G6740,G21754);
  nand GNAME5169(G5169,G7815,G1585);
  nand GNAME5170(G5170,G21627,G1582);
  nand GNAME5171(G5171,G21786,G4992);
  nand GNAME5172(G5172,G8263,G1584);
  nand GNAME5173(G5173,G6741,G7472);
  nand GNAME5174(G5174,G6740,G21755);
  nand GNAME5175(G5175,G7814,G1585);
  nand GNAME5176(G5176,G21628,G1582);
  nand GNAME5177(G5177,G21787,G4992);
  nand GNAME5178(G5178,G8209,G1584);
  nand GNAME5179(G5179,G6741,G7441);
  nand GNAME5180(G5180,G6740,G21756);
  nand GNAME5181(G5181,G7777,G1585);
  nand GNAME5182(G5182,G21629,G1582);
  nand GNAME5183(G5183,G21788,G4992);
  nand GNAME5184(G5184,G8210,G1584);
  nand GNAME5185(G5185,G6741,G7442);
  nand GNAME5186(G5186,G6740,G21757);
  nand GNAME5187(G5187,G7778,G1585);
  nand GNAME5188(G5188,G21630,G1582);
  nand GNAME5189(G5189,G21789,G4992);
  nor GNAME5190(G5190,G1206,G1207);
  or GNAME5191(G5191,G1542,G1587);
  nand GNAME5192(G5192,G1586,G21792);
  nand GNAME5193(G5193,G1257,G1506);
  or GNAME5194(G5194,G1502,G1545);
  nand GNAME5195(G5195,G5193,G21795);
  or GNAME5196(G5196,G2300,G1571);
  nand GNAME5197(G5197,G5196,G1283);
  nand GNAME5198(G5198,G5197,G1588);
  nand GNAME5199(G5199,G1283,G2297);
  nand GNAME5200(G5200,G5199,G1545);
  nand GNAME5201(G5201,G1502,G5200);
  nand GNAME5202(G5202,G1282,G5198);
  nand GNAME5203(G5203,G5201,G5202);
  nand GNAME5204(G5204,G1257,G5203);
  nand GNAME5205(G5205,G5193,G21796);
  nand GNAME5206(G5206,G1292,G1202,G21427);
  or GNAME5207(G5207,G21425,G1270);
  nand GNAME5208(G5208,G1248,G2545);
  nand GNAME5209(G5209,G5208,G2253);
  nand GNAME5210(G5210,G2545,G1276,G1248);
  nand GNAME5211(G5211,G1246,G5209);
  nand GNAME5212(G5212,G1202,G5210,G5211,G21426);
  nand GNAME5213(G5213,G5212,G21428);
  and GNAME5214(G5214,G5213,G2317);
  nand GNAME5215(G5215,G1256,G1506);
  nand GNAME5216(G5216,G5215,G21801);
  or GNAME5217(G5217,G1269,G1535);
  nand GNAME5218(G5218,G21392,G21802);
  nor GNAME5219(G5219,G1209,G1264,G682);
  nand GNAME5220(G5220,G21549,G1592);
  nand GNAME5221(G5221,G21541,G1594);
  nand GNAME5222(G5222,G21533,G1596);
  nand GNAME5223(G5223,G21525,G1597);
  nand GNAME5224(G5224,G21517,G1599);
  nand GNAME5225(G5225,G21509,G1601);
  nand GNAME5226(G5226,G21501,G1602);
  nand GNAME5227(G5227,G21493,G1603);
  nand GNAME5228(G5228,G21429,G1605);
  nand GNAME5229(G5229,G21437,G1606);
  nand GNAME5230(G5230,G21445,G1608);
  nand GNAME5231(G5231,G21453,G1609);
  nand GNAME5232(G5232,G21461,G1610);
  nand GNAME5233(G5233,G21469,G1611);
  nand GNAME5234(G5234,G21477,G1612);
  nand GNAME5235(G5235,G21485,G1613);
  nand GNAME5236(G5236,G21550,G1592);
  nand GNAME5237(G5237,G21542,G1594);
  nand GNAME5238(G5238,G21534,G1596);
  nand GNAME5239(G5239,G21526,G1597);
  nand GNAME5240(G5240,G21518,G1599);
  nand GNAME5241(G5241,G21510,G1601);
  nand GNAME5242(G5242,G21502,G1602);
  nand GNAME5243(G5243,G21494,G1603);
  nand GNAME5244(G5244,G21430,G1605);
  nand GNAME5245(G5245,G21438,G1606);
  nand GNAME5246(G5246,G21446,G1608);
  nand GNAME5247(G5247,G21454,G1609);
  nand GNAME5248(G5248,G21462,G1610);
  nand GNAME5249(G5249,G21470,G1611);
  nand GNAME5250(G5250,G21478,G1612);
  nand GNAME5251(G5251,G21486,G1613);
  nand GNAME5252(G5252,G21551,G1592);
  nand GNAME5253(G5253,G21543,G1594);
  nand GNAME5254(G5254,G21535,G1596);
  nand GNAME5255(G5255,G21527,G1597);
  nand GNAME5256(G5256,G21519,G1599);
  nand GNAME5257(G5257,G21511,G1601);
  nand GNAME5258(G5258,G21503,G1602);
  nand GNAME5259(G5259,G21495,G1603);
  nand GNAME5260(G5260,G21431,G1605);
  nand GNAME5261(G5261,G21439,G1606);
  nand GNAME5262(G5262,G21447,G1608);
  nand GNAME5263(G5263,G21455,G1609);
  nand GNAME5264(G5264,G21463,G1610);
  nand GNAME5265(G5265,G21471,G1611);
  nand GNAME5266(G5266,G21479,G1612);
  nand GNAME5267(G5267,G21487,G1613);
  nand GNAME5268(G5268,G21552,G1592);
  nand GNAME5269(G5269,G21544,G1594);
  nand GNAME5270(G5270,G21536,G1596);
  nand GNAME5271(G5271,G21528,G1597);
  nand GNAME5272(G5272,G21520,G1599);
  nand GNAME5273(G5273,G21512,G1601);
  nand GNAME5274(G5274,G21504,G1602);
  nand GNAME5275(G5275,G21496,G1603);
  nand GNAME5276(G5276,G21432,G1605);
  nand GNAME5277(G5277,G21440,G1606);
  nand GNAME5278(G5278,G21448,G1608);
  nand GNAME5279(G5279,G21456,G1609);
  nand GNAME5280(G5280,G21464,G1610);
  nand GNAME5281(G5281,G21472,G1611);
  nand GNAME5282(G5282,G21480,G1612);
  nand GNAME5283(G5283,G21488,G1613);
  nand GNAME5284(G5284,G21553,G1592);
  nand GNAME5285(G5285,G21545,G1594);
  nand GNAME5286(G5286,G21537,G1596);
  nand GNAME5287(G5287,G21529,G1597);
  nand GNAME5288(G5288,G21521,G1599);
  nand GNAME5289(G5289,G21513,G1601);
  nand GNAME5290(G5290,G21505,G1602);
  nand GNAME5291(G5291,G21497,G1603);
  nand GNAME5292(G5292,G21433,G1605);
  nand GNAME5293(G5293,G21441,G1606);
  nand GNAME5294(G5294,G21449,G1608);
  nand GNAME5295(G5295,G21457,G1609);
  nand GNAME5296(G5296,G21465,G1610);
  nand GNAME5297(G5297,G21473,G1611);
  nand GNAME5298(G5298,G21481,G1612);
  nand GNAME5299(G5299,G21489,G1613);
  nand GNAME5300(G5300,G21554,G1592);
  nand GNAME5301(G5301,G21546,G1594);
  nand GNAME5302(G5302,G21538,G1596);
  nand GNAME5303(G5303,G21530,G1597);
  nand GNAME5304(G5304,G21522,G1599);
  nand GNAME5305(G5305,G21514,G1601);
  nand GNAME5306(G5306,G21506,G1602);
  nand GNAME5307(G5307,G21498,G1603);
  nand GNAME5308(G5308,G21434,G1605);
  nand GNAME5309(G5309,G21442,G1606);
  nand GNAME5310(G5310,G21450,G1608);
  nand GNAME5311(G5311,G21458,G1609);
  nand GNAME5312(G5312,G21466,G1610);
  nand GNAME5313(G5313,G21474,G1611);
  nand GNAME5314(G5314,G21482,G1612);
  nand GNAME5315(G5315,G21490,G1613);
  nand GNAME5316(G5316,G21555,G1592);
  nand GNAME5317(G5317,G21547,G1594);
  nand GNAME5318(G5318,G21539,G1596);
  nand GNAME5319(G5319,G21531,G1597);
  nand GNAME5320(G5320,G21523,G1599);
  nand GNAME5321(G5321,G21515,G1601);
  nand GNAME5322(G5322,G21507,G1602);
  nand GNAME5323(G5323,G21499,G1603);
  nand GNAME5324(G5324,G21435,G1605);
  nand GNAME5325(G5325,G21443,G1606);
  nand GNAME5326(G5326,G21451,G1608);
  nand GNAME5327(G5327,G21459,G1609);
  nand GNAME5328(G5328,G21467,G1610);
  nand GNAME5329(G5329,G21475,G1611);
  nand GNAME5330(G5330,G21483,G1612);
  nand GNAME5331(G5331,G21491,G1613);
  nand GNAME5332(G5332,G21556,G1592);
  nand GNAME5333(G5333,G21548,G1594);
  nand GNAME5334(G5334,G21540,G1596);
  nand GNAME5335(G5335,G21532,G1597);
  nand GNAME5336(G5336,G21524,G1599);
  nand GNAME5337(G5337,G21516,G1601);
  nand GNAME5338(G5338,G21508,G1602);
  nand GNAME5339(G5339,G21500,G1603);
  nand GNAME5340(G5340,G21436,G1605);
  nand GNAME5341(G5341,G21444,G1606);
  nand GNAME5342(G5342,G21452,G1608);
  nand GNAME5343(G5343,G21460,G1609);
  nand GNAME5344(G5344,G21468,G1610);
  nand GNAME5345(G5345,G21476,G1611);
  nand GNAME5346(G5346,G21484,G1612);
  nand GNAME5347(G5347,G21492,G1613);
  nand GNAME5348(G5348,G21429,G1615);
  nand GNAME5349(G5349,G21437,G1616);
  nand GNAME5350(G5350,G21445,G1617);
  nand GNAME5351(G5351,G21453,G1618);
  nand GNAME5352(G5352,G21461,G1620);
  nand GNAME5353(G5353,G21469,G1621);
  nand GNAME5354(G5354,G21477,G1622);
  nand GNAME5355(G5355,G21485,G1623);
  nand GNAME5356(G5356,G21549,G1626);
  nand GNAME5357(G5357,G21541,G1627);
  nand GNAME5358(G5358,G21533,G1628);
  nand GNAME5359(G5359,G21525,G1629);
  nand GNAME5360(G5360,G21517,G1631);
  nand GNAME5361(G5361,G21509,G1632);
  nand GNAME5362(G5362,G21501,G1633);
  nand GNAME5363(G5363,G21493,G1634);
  nand GNAME5364(G5364,G21430,G1615);
  nand GNAME5365(G5365,G21438,G1616);
  nand GNAME5366(G5366,G21446,G1617);
  nand GNAME5367(G5367,G21454,G1618);
  nand GNAME5368(G5368,G21462,G1620);
  nand GNAME5369(G5369,G21470,G1621);
  nand GNAME5370(G5370,G21478,G1622);
  nand GNAME5371(G5371,G21486,G1623);
  nand GNAME5372(G5372,G21550,G1626);
  nand GNAME5373(G5373,G21542,G1627);
  nand GNAME5374(G5374,G21534,G1628);
  nand GNAME5375(G5375,G21526,G1629);
  nand GNAME5376(G5376,G21518,G1631);
  nand GNAME5377(G5377,G21510,G1632);
  nand GNAME5378(G5378,G21502,G1633);
  nand GNAME5379(G5379,G21494,G1634);
  nand GNAME5380(G5380,G21431,G1615);
  nand GNAME5381(G5381,G21439,G1616);
  nand GNAME5382(G5382,G21447,G1617);
  nand GNAME5383(G5383,G21455,G1618);
  nand GNAME5384(G5384,G21463,G1620);
  nand GNAME5385(G5385,G21471,G1621);
  nand GNAME5386(G5386,G21479,G1622);
  nand GNAME5387(G5387,G21487,G1623);
  nand GNAME5388(G5388,G21551,G1626);
  nand GNAME5389(G5389,G21543,G1627);
  nand GNAME5390(G5390,G21535,G1628);
  nand GNAME5391(G5391,G21527,G1629);
  nand GNAME5392(G5392,G21519,G1631);
  nand GNAME5393(G5393,G21511,G1632);
  nand GNAME5394(G5394,G21503,G1633);
  nand GNAME5395(G5395,G21495,G1634);
  nand GNAME5396(G5396,G21432,G1615);
  nand GNAME5397(G5397,G21440,G1616);
  nand GNAME5398(G5398,G21448,G1617);
  nand GNAME5399(G5399,G21456,G1618);
  nand GNAME5400(G5400,G21464,G1620);
  nand GNAME5401(G5401,G21472,G1621);
  nand GNAME5402(G5402,G21480,G1622);
  nand GNAME5403(G5403,G21488,G1623);
  nand GNAME5404(G5404,G21552,G1626);
  nand GNAME5405(G5405,G21544,G1627);
  nand GNAME5406(G5406,G21536,G1628);
  nand GNAME5407(G5407,G21528,G1629);
  nand GNAME5408(G5408,G21520,G1631);
  nand GNAME5409(G5409,G21512,G1632);
  nand GNAME5410(G5410,G21504,G1633);
  nand GNAME5411(G5411,G21496,G1634);
  nand GNAME5412(G5412,G21433,G1615);
  nand GNAME5413(G5413,G21441,G1616);
  nand GNAME5414(G5414,G21449,G1617);
  nand GNAME5415(G5415,G21457,G1618);
  nand GNAME5416(G5416,G21465,G1620);
  nand GNAME5417(G5417,G21473,G1621);
  nand GNAME5418(G5418,G21481,G1622);
  nand GNAME5419(G5419,G21489,G1623);
  nand GNAME5420(G5420,G21553,G1626);
  nand GNAME5421(G5421,G21545,G1627);
  nand GNAME5422(G5422,G21537,G1628);
  nand GNAME5423(G5423,G21529,G1629);
  nand GNAME5424(G5424,G21521,G1631);
  nand GNAME5425(G5425,G21513,G1632);
  nand GNAME5426(G5426,G21505,G1633);
  nand GNAME5427(G5427,G21497,G1634);
  nand GNAME5428(G5428,G21434,G1615);
  nand GNAME5429(G5429,G21442,G1616);
  nand GNAME5430(G5430,G21450,G1617);
  nand GNAME5431(G5431,G21458,G1618);
  nand GNAME5432(G5432,G21466,G1620);
  nand GNAME5433(G5433,G21474,G1621);
  nand GNAME5434(G5434,G21482,G1622);
  nand GNAME5435(G5435,G21490,G1623);
  nand GNAME5436(G5436,G21554,G1626);
  nand GNAME5437(G5437,G21546,G1627);
  nand GNAME5438(G5438,G21538,G1628);
  nand GNAME5439(G5439,G21530,G1629);
  nand GNAME5440(G5440,G21522,G1631);
  nand GNAME5441(G5441,G21514,G1632);
  nand GNAME5442(G5442,G21506,G1633);
  nand GNAME5443(G5443,G21498,G1634);
  nand GNAME5444(G5444,G21435,G1615);
  nand GNAME5445(G5445,G21443,G1616);
  nand GNAME5446(G5446,G21451,G1617);
  nand GNAME5447(G5447,G21459,G1618);
  nand GNAME5448(G5448,G21467,G1620);
  nand GNAME5449(G5449,G21475,G1621);
  nand GNAME5450(G5450,G21483,G1622);
  nand GNAME5451(G5451,G21491,G1623);
  nand GNAME5452(G5452,G21555,G1626);
  nand GNAME5453(G5453,G21547,G1627);
  nand GNAME5454(G5454,G21539,G1628);
  nand GNAME5455(G5455,G21531,G1629);
  nand GNAME5456(G5456,G21523,G1631);
  nand GNAME5457(G5457,G21515,G1632);
  nand GNAME5458(G5458,G21507,G1633);
  nand GNAME5459(G5459,G21499,G1634);
  nand GNAME5460(G5460,G21436,G1615);
  nand GNAME5461(G5461,G21444,G1616);
  nand GNAME5462(G5462,G21452,G1617);
  nand GNAME5463(G5463,G21460,G1618);
  nand GNAME5464(G5464,G21468,G1620);
  nand GNAME5465(G5465,G21476,G1621);
  nand GNAME5466(G5466,G21484,G1622);
  nand GNAME5467(G5467,G21492,G1623);
  nand GNAME5468(G5468,G21556,G1626);
  nand GNAME5469(G5469,G21548,G1627);
  nand GNAME5470(G5470,G21540,G1628);
  nand GNAME5471(G5471,G21532,G1629);
  nand GNAME5472(G5472,G21524,G1631);
  nand GNAME5473(G5473,G21516,G1632);
  nand GNAME5474(G5474,G21508,G1633);
  nand GNAME5475(G5475,G21500,G1634);
  nand GNAME5476(G5476,G21549,G1500);
  nand GNAME5477(G5477,G21541,G1492);
  nand GNAME5478(G5478,G21533,G1484);
  nand GNAME5479(G5479,G21525,G1476);
  nand GNAME5480(G5480,G21517,G1467);
  nand GNAME5481(G5481,G21509,G1459);
  nand GNAME5482(G5482,G21501,G1450);
  nand GNAME5483(G5483,G21493,G1442);
  nand GNAME5484(G5484,G21485,G1431);
  nand GNAME5485(G5485,G21477,G1421);
  nand GNAME5486(G5486,G21469,G1411);
  nand GNAME5487(G5487,G21461,G1400);
  nand GNAME5488(G5488,G21453,G1387);
  nand GNAME5489(G5489,G21445,G1376);
  nand GNAME5490(G5490,G21437,G1362);
  nand GNAME5491(G5491,G21429,G1326);
  nand GNAME5492(G5492,G2074,G2075,G2076,G2077);
  nand GNAME5493(G5493,G21550,G1500);
  nand GNAME5494(G5494,G21542,G1492);
  nand GNAME5495(G5495,G21534,G1484);
  nand GNAME5496(G5496,G21526,G1476);
  nand GNAME5497(G5497,G21518,G1467);
  nand GNAME5498(G5498,G21510,G1459);
  nand GNAME5499(G5499,G21502,G1450);
  nand GNAME5500(G5500,G21494,G1442);
  nand GNAME5501(G5501,G21486,G1431);
  nand GNAME5502(G5502,G21478,G1421);
  nand GNAME5503(G5503,G21470,G1411);
  nand GNAME5504(G5504,G21462,G1400);
  nand GNAME5505(G5505,G21454,G1387);
  nand GNAME5506(G5506,G21446,G1376);
  nand GNAME5507(G5507,G21438,G1362);
  nand GNAME5508(G5508,G21430,G1326);
  nand GNAME5509(G5509,G2078,G2079,G2080,G2081);
  nand GNAME5510(G5510,G21551,G1500);
  nand GNAME5511(G5511,G21543,G1492);
  nand GNAME5512(G5512,G21535,G1484);
  nand GNAME5513(G5513,G21527,G1476);
  nand GNAME5514(G5514,G21519,G1467);
  nand GNAME5515(G5515,G21511,G1459);
  nand GNAME5516(G5516,G21503,G1450);
  nand GNAME5517(G5517,G21495,G1442);
  nand GNAME5518(G5518,G21487,G1431);
  nand GNAME5519(G5519,G21479,G1421);
  nand GNAME5520(G5520,G21471,G1411);
  nand GNAME5521(G5521,G21463,G1400);
  nand GNAME5522(G5522,G21455,G1387);
  nand GNAME5523(G5523,G21447,G1376);
  nand GNAME5524(G5524,G21439,G1362);
  nand GNAME5525(G5525,G21431,G1326);
  nand GNAME5526(G5526,G2082,G2083,G2084,G2085);
  nand GNAME5527(G5527,G21552,G1500);
  nand GNAME5528(G5528,G21544,G1492);
  nand GNAME5529(G5529,G21536,G1484);
  nand GNAME5530(G5530,G21528,G1476);
  nand GNAME5531(G5531,G21520,G1467);
  nand GNAME5532(G5532,G21512,G1459);
  nand GNAME5533(G5533,G21504,G1450);
  nand GNAME5534(G5534,G21496,G1442);
  nand GNAME5535(G5535,G21488,G1431);
  nand GNAME5536(G5536,G21480,G1421);
  nand GNAME5537(G5537,G21472,G1411);
  nand GNAME5538(G5538,G21464,G1400);
  nand GNAME5539(G5539,G21456,G1387);
  nand GNAME5540(G5540,G21448,G1376);
  nand GNAME5541(G5541,G21440,G1362);
  nand GNAME5542(G5542,G21432,G1326);
  nand GNAME5543(G5543,G2086,G2087,G2088,G2089);
  nand GNAME5544(G5544,G21553,G1500);
  nand GNAME5545(G5545,G21545,G1492);
  nand GNAME5546(G5546,G21537,G1484);
  nand GNAME5547(G5547,G21529,G1476);
  nand GNAME5548(G5548,G21521,G1467);
  nand GNAME5549(G5549,G21513,G1459);
  nand GNAME5550(G5550,G21505,G1450);
  nand GNAME5551(G5551,G21497,G1442);
  nand GNAME5552(G5552,G21489,G1431);
  nand GNAME5553(G5553,G21481,G1421);
  nand GNAME5554(G5554,G21473,G1411);
  nand GNAME5555(G5555,G21465,G1400);
  nand GNAME5556(G5556,G21457,G1387);
  nand GNAME5557(G5557,G21449,G1376);
  nand GNAME5558(G5558,G21441,G1362);
  nand GNAME5559(G5559,G21433,G1326);
  nand GNAME5560(G5560,G2090,G2091,G2092,G2093);
  nand GNAME5561(G5561,G21554,G1500);
  nand GNAME5562(G5562,G21546,G1492);
  nand GNAME5563(G5563,G21538,G1484);
  nand GNAME5564(G5564,G21530,G1476);
  nand GNAME5565(G5565,G21522,G1467);
  nand GNAME5566(G5566,G21514,G1459);
  nand GNAME5567(G5567,G21506,G1450);
  nand GNAME5568(G5568,G21498,G1442);
  nand GNAME5569(G5569,G21490,G1431);
  nand GNAME5570(G5570,G21482,G1421);
  nand GNAME5571(G5571,G21474,G1411);
  nand GNAME5572(G5572,G21466,G1400);
  nand GNAME5573(G5573,G21458,G1387);
  nand GNAME5574(G5574,G21450,G1376);
  nand GNAME5575(G5575,G21442,G1362);
  nand GNAME5576(G5576,G21434,G1326);
  nand GNAME5577(G5577,G2094,G2095,G2096,G2097);
  nand GNAME5578(G5578,G21555,G1500);
  nand GNAME5579(G5579,G21547,G1492);
  nand GNAME5580(G5580,G21539,G1484);
  nand GNAME5581(G5581,G21531,G1476);
  nand GNAME5582(G5582,G21523,G1467);
  nand GNAME5583(G5583,G21515,G1459);
  nand GNAME5584(G5584,G21507,G1450);
  nand GNAME5585(G5585,G21499,G1442);
  nand GNAME5586(G5586,G21491,G1431);
  nand GNAME5587(G5587,G21483,G1421);
  nand GNAME5588(G5588,G21475,G1411);
  nand GNAME5589(G5589,G21467,G1400);
  nand GNAME5590(G5590,G21459,G1387);
  nand GNAME5591(G5591,G21451,G1376);
  nand GNAME5592(G5592,G21443,G1362);
  nand GNAME5593(G5593,G21435,G1326);
  nand GNAME5594(G5594,G2098,G2099,G2100,G2101);
  nand GNAME5595(G5595,G21556,G1500);
  nand GNAME5596(G5596,G21548,G1492);
  nand GNAME5597(G5597,G21540,G1484);
  nand GNAME5598(G5598,G21532,G1476);
  nand GNAME5599(G5599,G21524,G1467);
  nand GNAME5600(G5600,G21516,G1459);
  nand GNAME5601(G5601,G21508,G1450);
  nand GNAME5602(G5602,G21500,G1442);
  nand GNAME5603(G5603,G21492,G1431);
  nand GNAME5604(G5604,G21484,G1421);
  nand GNAME5605(G5605,G21476,G1411);
  nand GNAME5606(G5606,G21468,G1400);
  nand GNAME5607(G5607,G21460,G1387);
  nand GNAME5608(G5608,G21452,G1376);
  nand GNAME5609(G5609,G21444,G1362);
  nand GNAME5610(G5610,G21436,G1326);
  nand GNAME5611(G5611,G2102,G2103,G2104,G2105);
  nand GNAME5612(G5612,G21493,G1637);
  nand GNAME5613(G5613,G21501,G1639);
  nand GNAME5614(G5614,G21509,G1641);
  nand GNAME5615(G5615,G21517,G1642);
  nand GNAME5616(G5616,G21525,G1644);
  nand GNAME5617(G5617,G21533,G1646);
  nand GNAME5618(G5618,G21541,G1647);
  nand GNAME5619(G5619,G21549,G1648);
  nand GNAME5620(G5620,G21485,G1650);
  nand GNAME5621(G5621,G21477,G1651);
  nand GNAME5622(G5622,G21469,G1653);
  nand GNAME5623(G5623,G21461,G1654);
  nand GNAME5624(G5624,G21453,G1655);
  nand GNAME5625(G5625,G21445,G1656);
  nand GNAME5626(G5626,G21437,G1657);
  nand GNAME5627(G5627,G21429,G1658);
  nand GNAME5628(G5628,G2106,G2107,G2108,G2109);
  nand GNAME5629(G5629,G21494,G1637);
  nand GNAME5630(G5630,G21502,G1639);
  nand GNAME5631(G5631,G21510,G1641);
  nand GNAME5632(G5632,G21518,G1642);
  nand GNAME5633(G5633,G21526,G1644);
  nand GNAME5634(G5634,G21534,G1646);
  nand GNAME5635(G5635,G21542,G1647);
  nand GNAME5636(G5636,G21550,G1648);
  nand GNAME5637(G5637,G21486,G1650);
  nand GNAME5638(G5638,G21478,G1651);
  nand GNAME5639(G5639,G21470,G1653);
  nand GNAME5640(G5640,G21462,G1654);
  nand GNAME5641(G5641,G21454,G1655);
  nand GNAME5642(G5642,G21446,G1656);
  nand GNAME5643(G5643,G21438,G1657);
  nand GNAME5644(G5644,G21430,G1658);
  nand GNAME5645(G5645,G2110,G2111,G2112,G2113);
  nand GNAME5646(G5646,G21495,G1637);
  nand GNAME5647(G5647,G21503,G1639);
  nand GNAME5648(G5648,G21511,G1641);
  nand GNAME5649(G5649,G21519,G1642);
  nand GNAME5650(G5650,G21527,G1644);
  nand GNAME5651(G5651,G21535,G1646);
  nand GNAME5652(G5652,G21543,G1647);
  nand GNAME5653(G5653,G21551,G1648);
  nand GNAME5654(G5654,G21487,G1650);
  nand GNAME5655(G5655,G21479,G1651);
  nand GNAME5656(G5656,G21471,G1653);
  nand GNAME5657(G5657,G21463,G1654);
  nand GNAME5658(G5658,G21455,G1655);
  nand GNAME5659(G5659,G21447,G1656);
  nand GNAME5660(G5660,G21439,G1657);
  nand GNAME5661(G5661,G21431,G1658);
  nand GNAME5662(G5662,G2114,G2115,G2116,G2117);
  nand GNAME5663(G5663,G21496,G1637);
  nand GNAME5664(G5664,G21504,G1639);
  nand GNAME5665(G5665,G21512,G1641);
  nand GNAME5666(G5666,G21520,G1642);
  nand GNAME5667(G5667,G21528,G1644);
  nand GNAME5668(G5668,G21536,G1646);
  nand GNAME5669(G5669,G21544,G1647);
  nand GNAME5670(G5670,G21552,G1648);
  nand GNAME5671(G5671,G21488,G1650);
  nand GNAME5672(G5672,G21480,G1651);
  nand GNAME5673(G5673,G21472,G1653);
  nand GNAME5674(G5674,G21464,G1654);
  nand GNAME5675(G5675,G21456,G1655);
  nand GNAME5676(G5676,G21448,G1656);
  nand GNAME5677(G5677,G21440,G1657);
  nand GNAME5678(G5678,G21432,G1658);
  nand GNAME5679(G5679,G2118,G2119,G2120,G2121);
  nand GNAME5680(G5680,G21497,G1637);
  nand GNAME5681(G5681,G21505,G1639);
  nand GNAME5682(G5682,G21513,G1641);
  nand GNAME5683(G5683,G21521,G1642);
  nand GNAME5684(G5684,G21529,G1644);
  nand GNAME5685(G5685,G21537,G1646);
  nand GNAME5686(G5686,G21545,G1647);
  nand GNAME5687(G5687,G21553,G1648);
  nand GNAME5688(G5688,G21489,G1650);
  nand GNAME5689(G5689,G21481,G1651);
  nand GNAME5690(G5690,G21473,G1653);
  nand GNAME5691(G5691,G21465,G1654);
  nand GNAME5692(G5692,G21457,G1655);
  nand GNAME5693(G5693,G21449,G1656);
  nand GNAME5694(G5694,G21441,G1657);
  nand GNAME5695(G5695,G21433,G1658);
  nand GNAME5696(G5696,G2122,G2123,G2124,G2125);
  nand GNAME5697(G5697,G21498,G1637);
  nand GNAME5698(G5698,G21506,G1639);
  nand GNAME5699(G5699,G21514,G1641);
  nand GNAME5700(G5700,G21522,G1642);
  nand GNAME5701(G5701,G21530,G1644);
  nand GNAME5702(G5702,G21538,G1646);
  nand GNAME5703(G5703,G21546,G1647);
  nand GNAME5704(G5704,G21554,G1648);
  nand GNAME5705(G5705,G21490,G1650);
  nand GNAME5706(G5706,G21482,G1651);
  nand GNAME5707(G5707,G21474,G1653);
  nand GNAME5708(G5708,G21466,G1654);
  nand GNAME5709(G5709,G21458,G1655);
  nand GNAME5710(G5710,G21450,G1656);
  nand GNAME5711(G5711,G21442,G1657);
  nand GNAME5712(G5712,G21434,G1658);
  nand GNAME5713(G5713,G2126,G2127,G2128,G2129);
  nand GNAME5714(G5714,G21499,G1637);
  nand GNAME5715(G5715,G21507,G1639);
  nand GNAME5716(G5716,G21515,G1641);
  nand GNAME5717(G5717,G21523,G1642);
  nand GNAME5718(G5718,G21531,G1644);
  nand GNAME5719(G5719,G21539,G1646);
  nand GNAME5720(G5720,G21547,G1647);
  nand GNAME5721(G5721,G21555,G1648);
  nand GNAME5722(G5722,G21491,G1650);
  nand GNAME5723(G5723,G21483,G1651);
  nand GNAME5724(G5724,G21475,G1653);
  nand GNAME5725(G5725,G21467,G1654);
  nand GNAME5726(G5726,G21459,G1655);
  nand GNAME5727(G5727,G21451,G1656);
  nand GNAME5728(G5728,G21443,G1657);
  nand GNAME5729(G5729,G21435,G1658);
  nand GNAME5730(G5730,G2130,G2131,G2132,G2133);
  nand GNAME5731(G5731,G21500,G1637);
  nand GNAME5732(G5732,G21508,G1639);
  nand GNAME5733(G5733,G21516,G1641);
  nand GNAME5734(G5734,G21524,G1642);
  nand GNAME5735(G5735,G21532,G1644);
  nand GNAME5736(G5736,G21540,G1646);
  nand GNAME5737(G5737,G21548,G1647);
  nand GNAME5738(G5738,G21556,G1648);
  nand GNAME5739(G5739,G21492,G1650);
  nand GNAME5740(G5740,G21484,G1651);
  nand GNAME5741(G5741,G21476,G1653);
  nand GNAME5742(G5742,G21468,G1654);
  nand GNAME5743(G5743,G21460,G1655);
  nand GNAME5744(G5744,G21452,G1656);
  nand GNAME5745(G5745,G21444,G1657);
  nand GNAME5746(G5746,G21436,G1658);
  nand GNAME5747(G5747,G2134,G2135,G2136,G2137);
  nand GNAME5748(G5748,G2312,G2310,G2311);
  or GNAME5749(G5749,G1662,G1687);
  nand GNAME5750(G5750,G5749,G7810);
  nand GNAME5751(G5751,G5748,G21576);
  nand GNAME5752(G5752,G1260,G8539);
  nand GNAME5753(G5753,G21767,G1660);
  nand GNAME5754(G5754,G7468,G1661);
  nand GNAME5755(G5755,G5749,G7811);
  nand GNAME5756(G5756,G5748,G21575);
  nand GNAME5757(G5757,G1260,G8579);
  nand GNAME5758(G5758,G21766,G1660);
  nand GNAME5759(G5759,G7469,G1661);
  nand GNAME5760(G5760,G5749,G7781);
  nand GNAME5761(G5761,G5748,G21574);
  nand GNAME5762(G5762,G1260,G7781);
  nand GNAME5763(G5763,G21765,G1660);
  nand GNAME5764(G5764,G7445,G1661);
  nand GNAME5765(G5765,G5749,G7780);
  nand GNAME5766(G5766,G5748,G21573);
  nand GNAME5767(G5767,G1260,G7780);
  nand GNAME5768(G5768,G21764,G1660);
  nand GNAME5769(G5769,G7444,G1661);
  nand GNAME5770(G5770,G5749,G7812);
  nand GNAME5771(G5771,G5748,G21572);
  nand GNAME5772(G5772,G1260,G7812);
  nand GNAME5773(G5773,G21763,G1660);
  nand GNAME5774(G5774,G7470,G1661);
  nand GNAME5775(G5775,G5749,G7813);
  nand GNAME5776(G5776,G5748,G21571);
  nand GNAME5777(G5777,G1260,G7813);
  nand GNAME5778(G5778,G21762,G1660);
  nand GNAME5779(G5779,G7471,G1661);
  nand GNAME5780(G5780,G5749,G7778);
  nand GNAME5781(G5781,G5748,G21598);
  nand GNAME5782(G5782,G21789,G1660);
  nand GNAME5783(G5783,G7442,G1661);
  nand GNAME5784(G5784,G5749,G7777);
  nand GNAME5785(G5785,G5748,G21597);
  nand GNAME5786(G5786,G1260,G8580);
  nand GNAME5787(G5787,G21788,G1660);
  nand GNAME5788(G5788,G7441,G1661);
  nand GNAME5789(G5789,G5749,G7779);
  nand GNAME5790(G5790,G5748,G21570);
  nand GNAME5791(G5791,G1260,G7779);
  nand GNAME5792(G5792,G21761,G1660);
  nand GNAME5793(G5793,G7443,G1661);
  nand GNAME5794(G5794,G5749,G7814);
  nand GNAME5795(G5795,G5748,G21596);
  nand GNAME5796(G5796,G1260,G8581);
  nand GNAME5797(G5797,G21787,G1660);
  nand GNAME5798(G5798,G7472,G1661);
  nand GNAME5799(G5799,G5749,G7815);
  nand GNAME5800(G5800,G5748,G21595);
  nand GNAME5801(G5801,G1260,G8582);
  nand GNAME5802(G5802,G21786,G1660);
  nand GNAME5803(G5803,G7473,G1661);
  nand GNAME5804(G5804,G5749,G7816);
  nand GNAME5805(G5805,G5748,G21594);
  nand GNAME5806(G5806,G1260,G8583);
  nand GNAME5807(G5807,G21785,G1660);
  nand GNAME5808(G5808,G7474,G1661);
  nand GNAME5809(G5809,G5749,G7817);
  nand GNAME5810(G5810,G5748,G21593);
  nand GNAME5811(G5811,G1260,G8584);
  nand GNAME5812(G5812,G21784,G1660);
  nand GNAME5813(G5813,G7475,G1661);
  nand GNAME5814(G5814,G5749,G7818);
  nand GNAME5815(G5815,G5748,G21592);
  nand GNAME5816(G5816,G1260,G8585);
  nand GNAME5817(G5817,G21783,G1660);
  nand GNAME5818(G5818,G7476,G1661);
  nand GNAME5819(G5819,G5749,G7819);
  nand GNAME5820(G5820,G5748,G21591);
  nand GNAME5821(G5821,G1260,G8586);
  nand GNAME5822(G5822,G21782,G1660);
  nand GNAME5823(G5823,G7477,G1661);
  nand GNAME5824(G5824,G5749,G7820);
  nand GNAME5825(G5825,G5748,G21590);
  nand GNAME5826(G5826,G1260,G8587);
  nand GNAME5827(G5827,G21781,G1660);
  nand GNAME5828(G5828,G7478,G1661);
  nand GNAME5829(G5829,G5749,G7821);
  nand GNAME5830(G5830,G5748,G21589);
  nand GNAME5831(G5831,G1260,G8588);
  nand GNAME5832(G5832,G21780,G1660);
  nand GNAME5833(G5833,G7479,G1661);
  nand GNAME5834(G5834,G5749,G7822);
  nand GNAME5835(G5835,G5748,G21588);
  nand GNAME5836(G5836,G1260,G8589);
  nand GNAME5837(G5837,G21779,G1660);
  nand GNAME5838(G5838,G7480,G1661);
  nand GNAME5839(G5839,G5749,G7823);
  nand GNAME5840(G5840,G5748,G21587);
  nand GNAME5841(G5841,G1260,G8590);
  nand GNAME5842(G5842,G21778,G1660);
  nand GNAME5843(G5843,G7481,G1661);
  nand GNAME5844(G5844,G5749,G7776);
  nand GNAME5845(G5845,G5748,G21569);
  nand GNAME5846(G5846,G1260,G7776);
  nand GNAME5847(G5847,G21760,G1660);
  nand GNAME5848(G5848,G7440,G1661);
  nand GNAME5849(G5849,G5749,G7825);
  nand GNAME5850(G5850,G5748,G21586);
  nand GNAME5851(G5851,G1260,G8591);
  nand GNAME5852(G5852,G21777,G1660);
  nand GNAME5853(G5853,G7483,G1661);
  nand GNAME5854(G5854,G5749,G7826);
  nand GNAME5855(G5855,G5748,G21585);
  nand GNAME5856(G5856,G1260,G8592);
  nand GNAME5857(G5857,G21776,G1660);
  nand GNAME5858(G5858,G7484,G1661);
  nand GNAME5859(G5859,G5749,G7827);
  nand GNAME5860(G5860,G5748,G21584);
  nand GNAME5861(G5861,G1260,G8593);
  nand GNAME5862(G5862,G21775,G1660);
  nand GNAME5863(G5863,G7485,G1661);
  nand GNAME5864(G5864,G5749,G7828);
  nand GNAME5865(G5865,G5748,G21583);
  nand GNAME5866(G5866,G1260,G8604);
  nand GNAME5867(G5867,G21774,G1660);
  nand GNAME5868(G5868,G7486,G1661);
  nand GNAME5869(G5869,G5749,G7829);
  nand GNAME5870(G5870,G5748,G21582);
  nand GNAME5871(G5871,G1260,G8538);
  nand GNAME5872(G5872,G21773,G1660);
  nand GNAME5873(G5873,G7487,G1661);
  nand GNAME5874(G5874,G5749,G7775);
  nand GNAME5875(G5875,G5748,G21581);
  nand GNAME5876(G5876,G1260,G8594);
  nand GNAME5877(G5877,G21772,G1660);
  nand GNAME5878(G5878,G7439,G1661);
  nand GNAME5879(G5879,G5749,G7830);
  nand GNAME5880(G5880,G5748,G21580);
  nand GNAME5881(G5881,G1260,G8595);
  nand GNAME5882(G5882,G21771,G1660);
  nand GNAME5883(G5883,G7488,G1661);
  nand GNAME5884(G5884,G5749,G7831);
  nand GNAME5885(G5885,G5748,G21579);
  nand GNAME5886(G5886,G1260,G8596);
  nand GNAME5887(G5887,G21770,G1660);
  nand GNAME5888(G5888,G7489,G1661);
  nand GNAME5889(G5889,G5749,G7774);
  nand GNAME5890(G5890,G5748,G21578);
  nand GNAME5891(G5891,G1260,G8597);
  nand GNAME5892(G5892,G21769,G1660);
  nand GNAME5893(G5893,G7438,G1661);
  nand GNAME5894(G5894,G5749,G7773);
  nand GNAME5895(G5895,G5748,G21577);
  nand GNAME5896(G5896,G1260,G8598);
  nand GNAME5897(G5897,G21768,G1660);
  nand GNAME5898(G5898,G7437,G1661);
  nand GNAME5899(G5899,G5749,G7824);
  nand GNAME5900(G5900,G5748,G21568);
  nand GNAME5901(G5901,G1260,G7824);
  nand GNAME5902(G5902,G21759,G1660);
  nand GNAME5903(G5903,G7482,G1661);
  nand GNAME5904(G5904,G5749,G7809);
  nand GNAME5905(G5905,G5748,G21567);
  nand GNAME5906(G5906,G1260,G7809);
  nand GNAME5907(G5907,G21758,G1660);
  nand GNAME5908(G5908,G7467,G1661);
  nand GNAME5909(G5909,G21549,G1691);
  nand GNAME5910(G5910,G21541,G1693);
  nand GNAME5911(G5911,G21533,G1695);
  nand GNAME5912(G5912,G21525,G1696);
  nand GNAME5913(G5913,G21517,G1698);
  nand GNAME5914(G5914,G21509,G1700);
  nand GNAME5915(G5915,G21501,G1701);
  nand GNAME5916(G5916,G21493,G1702);
  nand GNAME5917(G5917,G21485,G1704);
  nand GNAME5918(G5918,G21477,G1705);
  nand GNAME5919(G5919,G21469,G1707);
  nand GNAME5920(G5920,G21461,G1708);
  nand GNAME5921(G5921,G21453,G1709);
  nand GNAME5922(G5922,G21445,G1710);
  nand GNAME5923(G5923,G21437,G1711);
  nand GNAME5924(G5924,G21429,G1712);
  nand GNAME5925(G5925,G2147,G2148,G2149,G2150);
  nand GNAME5926(G5926,G21429,G2286);
  nand GNAME5927(G5927,G21437,G2285);
  nand GNAME5928(G5928,G21445,G2284);
  nand GNAME5929(G5929,G21453,G2283);
  nand GNAME5930(G5930,G21461,G2282);
  nand GNAME5931(G5931,G21469,G2281);
  nand GNAME5932(G5932,G21477,G2280);
  nand GNAME5933(G5933,G21485,G2279);
  nand GNAME5934(G5934,G21493,G2276);
  nand GNAME5935(G5935,G21501,G2275);
  nand GNAME5936(G5936,G21509,G2274);
  nand GNAME5937(G5937,G21517,G2273);
  nand GNAME5938(G5938,G21525,G2272);
  nand GNAME5939(G5939,G21533,G2271);
  nand GNAME5940(G5940,G21541,G2270);
  nand GNAME5941(G5941,G21549,G2269);
  nand GNAME5942(G5942,G2139,G2140,G2141,G2142);
  nand GNAME5943(G5943,G21429,G1665);
  nand GNAME5944(G5944,G21437,G1667);
  nand GNAME5945(G5945,G21445,G1669);
  nand GNAME5946(G5946,G21453,G1670);
  nand GNAME5947(G5947,G21461,G1672);
  nand GNAME5948(G5948,G21469,G1674);
  nand GNAME5949(G5949,G21477,G1675);
  nand GNAME5950(G5950,G21485,G1676);
  nand GNAME5951(G5951,G21493,G1678);
  nand GNAME5952(G5952,G21501,G1679);
  nand GNAME5953(G5953,G21509,G1681);
  nand GNAME5954(G5954,G21517,G1682);
  nand GNAME5955(G5955,G21525,G1683);
  nand GNAME5956(G5956,G21533,G1684);
  nand GNAME5957(G5957,G21541,G1685);
  nand GNAME5958(G5958,G21549,G1686);
  nand GNAME5959(G5959,G2143,G2144,G2145,G2146);
  nand GNAME5960(G5960,G1661,G7715);
  nand GNAME5961(G5961,G5942,G1662);
  nand GNAME5962(G5962,G5959,G1687);
  nand GNAME5963(G5963,G5925,G1260);
  nand GNAME5964(G5964,G21550,G1691);
  nand GNAME5965(G5965,G21542,G1693);
  nand GNAME5966(G5966,G21534,G1695);
  nand GNAME5967(G5967,G21526,G1696);
  nand GNAME5968(G5968,G21518,G1698);
  nand GNAME5969(G5969,G21510,G1700);
  nand GNAME5970(G5970,G21502,G1701);
  nand GNAME5971(G5971,G21494,G1702);
  nand GNAME5972(G5972,G21486,G1704);
  nand GNAME5973(G5973,G21478,G1705);
  nand GNAME5974(G5974,G21470,G1707);
  nand GNAME5975(G5975,G21462,G1708);
  nand GNAME5976(G5976,G21454,G1709);
  nand GNAME5977(G5977,G21446,G1710);
  nand GNAME5978(G5978,G21438,G1711);
  nand GNAME5979(G5979,G21430,G1712);
  nand GNAME5980(G5980,G2159,G2160,G2161,G2162);
  nand GNAME5981(G5981,G21430,G2286);
  nand GNAME5982(G5982,G21438,G2285);
  nand GNAME5983(G5983,G21446,G2284);
  nand GNAME5984(G5984,G21454,G2283);
  nand GNAME5985(G5985,G21462,G2282);
  nand GNAME5986(G5986,G21470,G2281);
  nand GNAME5987(G5987,G21478,G2280);
  nand GNAME5988(G5988,G21486,G2279);
  nand GNAME5989(G5989,G21494,G2276);
  nand GNAME5990(G5990,G21502,G2275);
  nand GNAME5991(G5991,G21510,G2274);
  nand GNAME5992(G5992,G21518,G2273);
  nand GNAME5993(G5993,G21526,G2272);
  nand GNAME5994(G5994,G21534,G2271);
  nand GNAME5995(G5995,G21542,G2270);
  nand GNAME5996(G5996,G21550,G2269);
  nand GNAME5997(G5997,G2151,G2152,G2153,G2154);
  nand GNAME5998(G5998,G21430,G1665);
  nand GNAME5999(G5999,G21438,G1667);
  nand GNAME6000(G6000,G21446,G1669);
  nand GNAME6001(G6001,G21454,G1670);
  nand GNAME6002(G6002,G21462,G1672);
  nand GNAME6003(G6003,G21470,G1674);
  nand GNAME6004(G6004,G21478,G1675);
  nand GNAME6005(G6005,G21486,G1676);
  nand GNAME6006(G6006,G21494,G1678);
  nand GNAME6007(G6007,G21502,G1679);
  nand GNAME6008(G6008,G21510,G1681);
  nand GNAME6009(G6009,G21518,G1682);
  nand GNAME6010(G6010,G21526,G1683);
  nand GNAME6011(G6011,G21534,G1684);
  nand GNAME6012(G6012,G21542,G1685);
  nand GNAME6013(G6013,G21550,G1686);
  nand GNAME6014(G6014,G2155,G2156,G2157,G2158);
  nand GNAME6015(G6015,G1661,G7713);
  nand GNAME6016(G6016,G5997,G1662);
  nand GNAME6017(G6017,G6014,G1687);
  nand GNAME6018(G6018,G5980,G1260);
  nand GNAME6019(G6019,G21551,G1691);
  nand GNAME6020(G6020,G21543,G1693);
  nand GNAME6021(G6021,G21535,G1695);
  nand GNAME6022(G6022,G21527,G1696);
  nand GNAME6023(G6023,G21519,G1698);
  nand GNAME6024(G6024,G21511,G1700);
  nand GNAME6025(G6025,G21503,G1701);
  nand GNAME6026(G6026,G21495,G1702);
  nand GNAME6027(G6027,G21487,G1704);
  nand GNAME6028(G6028,G21479,G1705);
  nand GNAME6029(G6029,G21471,G1707);
  nand GNAME6030(G6030,G21463,G1708);
  nand GNAME6031(G6031,G21455,G1709);
  nand GNAME6032(G6032,G21447,G1710);
  nand GNAME6033(G6033,G21439,G1711);
  nand GNAME6034(G6034,G21431,G1712);
  nand GNAME6035(G6035,G2171,G2172,G2173,G2174);
  nand GNAME6036(G6036,G21431,G2286);
  nand GNAME6037(G6037,G21439,G2285);
  nand GNAME6038(G6038,G21447,G2284);
  nand GNAME6039(G6039,G21455,G2283);
  nand GNAME6040(G6040,G21463,G2282);
  nand GNAME6041(G6041,G21471,G2281);
  nand GNAME6042(G6042,G21479,G2280);
  nand GNAME6043(G6043,G21487,G2279);
  nand GNAME6044(G6044,G21495,G2276);
  nand GNAME6045(G6045,G21503,G2275);
  nand GNAME6046(G6046,G21511,G2274);
  nand GNAME6047(G6047,G21519,G2273);
  nand GNAME6048(G6048,G21527,G2272);
  nand GNAME6049(G6049,G21535,G2271);
  nand GNAME6050(G6050,G21543,G2270);
  nand GNAME6051(G6051,G21551,G2269);
  nand GNAME6052(G6052,G2163,G2164,G2165,G2166);
  nand GNAME6053(G6053,G21431,G1665);
  nand GNAME6054(G6054,G21439,G1667);
  nand GNAME6055(G6055,G21447,G1669);
  nand GNAME6056(G6056,G21455,G1670);
  nand GNAME6057(G6057,G21463,G1672);
  nand GNAME6058(G6058,G21471,G1674);
  nand GNAME6059(G6059,G21479,G1675);
  nand GNAME6060(G6060,G21487,G1676);
  nand GNAME6061(G6061,G21495,G1678);
  nand GNAME6062(G6062,G21503,G1679);
  nand GNAME6063(G6063,G21511,G1681);
  nand GNAME6064(G6064,G21519,G1682);
  nand GNAME6065(G6065,G21527,G1683);
  nand GNAME6066(G6066,G21535,G1684);
  nand GNAME6067(G6067,G21543,G1685);
  nand GNAME6068(G6068,G21551,G1686);
  nand GNAME6069(G6069,G2167,G2168,G2169,G2170);
  nand GNAME6070(G6070,G1661,G7716);
  nand GNAME6071(G6071,G6052,G1662);
  nand GNAME6072(G6072,G6069,G1687);
  nand GNAME6073(G6073,G6035,G1260);
  nand GNAME6074(G6074,G21552,G1691);
  nand GNAME6075(G6075,G21544,G1693);
  nand GNAME6076(G6076,G21536,G1695);
  nand GNAME6077(G6077,G21528,G1696);
  nand GNAME6078(G6078,G21520,G1698);
  nand GNAME6079(G6079,G21512,G1700);
  nand GNAME6080(G6080,G21504,G1701);
  nand GNAME6081(G6081,G21496,G1702);
  nand GNAME6082(G6082,G21488,G1704);
  nand GNAME6083(G6083,G21480,G1705);
  nand GNAME6084(G6084,G21472,G1707);
  nand GNAME6085(G6085,G21464,G1708);
  nand GNAME6086(G6086,G21456,G1709);
  nand GNAME6087(G6087,G21448,G1710);
  nand GNAME6088(G6088,G21440,G1711);
  nand GNAME6089(G6089,G21432,G1712);
  nand GNAME6090(G6090,G2183,G2184,G2185,G2186);
  nand GNAME6091(G6091,G21432,G2286);
  nand GNAME6092(G6092,G21440,G2285);
  nand GNAME6093(G6093,G21448,G2284);
  nand GNAME6094(G6094,G21456,G2283);
  nand GNAME6095(G6095,G21464,G2282);
  nand GNAME6096(G6096,G21472,G2281);
  nand GNAME6097(G6097,G21480,G2280);
  nand GNAME6098(G6098,G21488,G2279);
  nand GNAME6099(G6099,G21496,G2276);
  nand GNAME6100(G6100,G21504,G2275);
  nand GNAME6101(G6101,G21512,G2274);
  nand GNAME6102(G6102,G21520,G2273);
  nand GNAME6103(G6103,G21528,G2272);
  nand GNAME6104(G6104,G21536,G2271);
  nand GNAME6105(G6105,G21544,G2270);
  nand GNAME6106(G6106,G21552,G2269);
  nand GNAME6107(G6107,G2175,G2176,G2177,G2178);
  nand GNAME6108(G6108,G21432,G1665);
  nand GNAME6109(G6109,G21440,G1667);
  nand GNAME6110(G6110,G21448,G1669);
  nand GNAME6111(G6111,G21456,G1670);
  nand GNAME6112(G6112,G21464,G1672);
  nand GNAME6113(G6113,G21472,G1674);
  nand GNAME6114(G6114,G21480,G1675);
  nand GNAME6115(G6115,G21488,G1676);
  nand GNAME6116(G6116,G21496,G1678);
  nand GNAME6117(G6117,G21504,G1679);
  nand GNAME6118(G6118,G21512,G1681);
  nand GNAME6119(G6119,G21520,G1682);
  nand GNAME6120(G6120,G21528,G1683);
  nand GNAME6121(G6121,G21536,G1684);
  nand GNAME6122(G6122,G21544,G1685);
  nand GNAME6123(G6123,G21552,G1686);
  nand GNAME6124(G6124,G2179,G2180,G2181,G2182);
  or GNAME6125(G6125,G2596,G7289);
  nand GNAME6126(G6126,G1661,G7720);
  nand GNAME6127(G6127,G6107,G1662);
  nand GNAME6128(G6128,G6124,G1687);
  nand GNAME6129(G6129,G6090,G1260);
  nand GNAME6130(G6130,G21553,G1691);
  nand GNAME6131(G6131,G21545,G1693);
  nand GNAME6132(G6132,G21537,G1695);
  nand GNAME6133(G6133,G21529,G1696);
  nand GNAME6134(G6134,G21521,G1698);
  nand GNAME6135(G6135,G21513,G1700);
  nand GNAME6136(G6136,G21505,G1701);
  nand GNAME6137(G6137,G21497,G1702);
  nand GNAME6138(G6138,G21489,G1704);
  nand GNAME6139(G6139,G21481,G1705);
  nand GNAME6140(G6140,G21473,G1707);
  nand GNAME6141(G6141,G21465,G1708);
  nand GNAME6142(G6142,G21457,G1709);
  nand GNAME6143(G6143,G21449,G1710);
  nand GNAME6144(G6144,G21441,G1711);
  nand GNAME6145(G6145,G21433,G1712);
  nand GNAME6146(G6146,G2195,G2196,G2197,G2198);
  nand GNAME6147(G6147,G21433,G2286);
  nand GNAME6148(G6148,G21441,G2285);
  nand GNAME6149(G6149,G21449,G2284);
  nand GNAME6150(G6150,G21457,G2283);
  nand GNAME6151(G6151,G21465,G2282);
  nand GNAME6152(G6152,G21473,G2281);
  nand GNAME6153(G6153,G21481,G2280);
  nand GNAME6154(G6154,G21489,G2279);
  nand GNAME6155(G6155,G21497,G2276);
  nand GNAME6156(G6156,G21505,G2275);
  nand GNAME6157(G6157,G21513,G2274);
  nand GNAME6158(G6158,G21521,G2273);
  nand GNAME6159(G6159,G21529,G2272);
  nand GNAME6160(G6160,G21537,G2271);
  nand GNAME6161(G6161,G21545,G2270);
  nand GNAME6162(G6162,G21553,G2269);
  nand GNAME6163(G6163,G2187,G2188,G2189,G2190);
  nand GNAME6164(G6164,G21433,G1665);
  nand GNAME6165(G6165,G21441,G1667);
  nand GNAME6166(G6166,G21449,G1669);
  nand GNAME6167(G6167,G21457,G1670);
  nand GNAME6168(G6168,G21465,G1672);
  nand GNAME6169(G6169,G21473,G1674);
  nand GNAME6170(G6170,G21481,G1675);
  nand GNAME6171(G6171,G21489,G1676);
  nand GNAME6172(G6172,G21497,G1678);
  nand GNAME6173(G6173,G21505,G1679);
  nand GNAME6174(G6174,G21513,G1681);
  nand GNAME6175(G6175,G21521,G1682);
  nand GNAME6176(G6176,G21529,G1683);
  nand GNAME6177(G6177,G21537,G1684);
  nand GNAME6178(G6178,G21545,G1685);
  nand GNAME6179(G6179,G21553,G1686);
  nand GNAME6180(G6180,G2191,G2192,G2193,G2194);
  nand GNAME6181(G6181,G1240,G21558);
  nand GNAME6182(G6182,G1661,G7718);
  nand GNAME6183(G6183,G6163,G1662);
  nand GNAME6184(G6184,G6180,G1687);
  nand GNAME6185(G6185,G6146,G1260);
  nand GNAME6186(G6186,G21554,G1691);
  nand GNAME6187(G6187,G21546,G1693);
  nand GNAME6188(G6188,G21538,G1695);
  nand GNAME6189(G6189,G21530,G1696);
  nand GNAME6190(G6190,G21522,G1698);
  nand GNAME6191(G6191,G21514,G1700);
  nand GNAME6192(G6192,G21506,G1701);
  nand GNAME6193(G6193,G21498,G1702);
  nand GNAME6194(G6194,G21490,G1704);
  nand GNAME6195(G6195,G21482,G1705);
  nand GNAME6196(G6196,G21474,G1707);
  nand GNAME6197(G6197,G21466,G1708);
  nand GNAME6198(G6198,G21458,G1709);
  nand GNAME6199(G6199,G21450,G1710);
  nand GNAME6200(G6200,G21442,G1711);
  nand GNAME6201(G6201,G21434,G1712);
  nand GNAME6202(G6202,G2207,G2208,G2209,G2210);
  nand GNAME6203(G6203,G21434,G2286);
  nand GNAME6204(G6204,G21442,G2285);
  nand GNAME6205(G6205,G21450,G2284);
  nand GNAME6206(G6206,G21458,G2283);
  nand GNAME6207(G6207,G21466,G2282);
  nand GNAME6208(G6208,G21474,G2281);
  nand GNAME6209(G6209,G21482,G2280);
  nand GNAME6210(G6210,G21490,G2279);
  nand GNAME6211(G6211,G21498,G2276);
  nand GNAME6212(G6212,G21506,G2275);
  nand GNAME6213(G6213,G21514,G2274);
  nand GNAME6214(G6214,G21522,G2273);
  nand GNAME6215(G6215,G21530,G2272);
  nand GNAME6216(G6216,G21538,G2271);
  nand GNAME6217(G6217,G21546,G2270);
  nand GNAME6218(G6218,G21554,G2269);
  nand GNAME6219(G6219,G2199,G2200,G2201,G2202);
  nand GNAME6220(G6220,G21434,G1665);
  nand GNAME6221(G6221,G21442,G1667);
  nand GNAME6222(G6222,G21450,G1669);
  nand GNAME6223(G6223,G21458,G1670);
  nand GNAME6224(G6224,G21466,G1672);
  nand GNAME6225(G6225,G21474,G1674);
  nand GNAME6226(G6226,G21482,G1675);
  nand GNAME6227(G6227,G21490,G1676);
  nand GNAME6228(G6228,G21498,G1678);
  nand GNAME6229(G6229,G21506,G1679);
  nand GNAME6230(G6230,G21514,G1681);
  nand GNAME6231(G6231,G21522,G1682);
  nand GNAME6232(G6232,G21530,G1683);
  nand GNAME6233(G6233,G21538,G1684);
  nand GNAME6234(G6234,G21546,G1685);
  nand GNAME6235(G6235,G21554,G1686);
  nand GNAME6236(G6236,G2203,G2204,G2205,G2206);
  nand GNAME6237(G6237,G1240,G21559);
  nand GNAME6238(G6238,G1661,G7719);
  nand GNAME6239(G6239,G6219,G1662);
  nand GNAME6240(G6240,G6236,G1687);
  nand GNAME6241(G6241,G6202,G1260);
  nand GNAME6242(G6242,G21555,G1691);
  nand GNAME6243(G6243,G21547,G1693);
  nand GNAME6244(G6244,G21539,G1695);
  nand GNAME6245(G6245,G21531,G1696);
  nand GNAME6246(G6246,G21523,G1698);
  nand GNAME6247(G6247,G21515,G1700);
  nand GNAME6248(G6248,G21507,G1701);
  nand GNAME6249(G6249,G21499,G1702);
  nand GNAME6250(G6250,G21491,G1704);
  nand GNAME6251(G6251,G21483,G1705);
  nand GNAME6252(G6252,G21475,G1707);
  nand GNAME6253(G6253,G21467,G1708);
  nand GNAME6254(G6254,G21459,G1709);
  nand GNAME6255(G6255,G21451,G1710);
  nand GNAME6256(G6256,G21443,G1711);
  nand GNAME6257(G6257,G21435,G1712);
  nand GNAME6258(G6258,G2220,G2221,G2222,G2223);
  nand GNAME6259(G6259,G21435,G2286);
  nand GNAME6260(G6260,G21443,G2285);
  nand GNAME6261(G6261,G21451,G2284);
  nand GNAME6262(G6262,G21459,G2283);
  nand GNAME6263(G6263,G21467,G2282);
  nand GNAME6264(G6264,G21475,G2281);
  nand GNAME6265(G6265,G21483,G2280);
  nand GNAME6266(G6266,G21491,G2279);
  nand GNAME6267(G6267,G21499,G2276);
  nand GNAME6268(G6268,G21507,G2275);
  nand GNAME6269(G6269,G21515,G2274);
  nand GNAME6270(G6270,G21523,G2273);
  nand GNAME6271(G6271,G21531,G2272);
  nand GNAME6272(G6272,G21539,G2271);
  nand GNAME6273(G6273,G21547,G2270);
  nand GNAME6274(G6274,G21555,G2269);
  nand GNAME6275(G6275,G2212,G2213,G2214,G2215);
  nand GNAME6276(G6276,G21435,G1665);
  nand GNAME6277(G6277,G21443,G1667);
  nand GNAME6278(G6278,G21451,G1669);
  nand GNAME6279(G6279,G21459,G1670);
  nand GNAME6280(G6280,G21467,G1672);
  nand GNAME6281(G6281,G21475,G1674);
  nand GNAME6282(G6282,G21483,G1675);
  nand GNAME6283(G6283,G21491,G1676);
  nand GNAME6284(G6284,G21499,G1678);
  nand GNAME6285(G6285,G21507,G1679);
  nand GNAME6286(G6286,G21515,G1681);
  nand GNAME6287(G6287,G21523,G1682);
  nand GNAME6288(G6288,G21531,G1683);
  nand GNAME6289(G6289,G21539,G1684);
  nand GNAME6290(G6290,G21547,G1685);
  nand GNAME6291(G6291,G21555,G1686);
  nand GNAME6292(G6292,G2216,G2217,G2218,G2219);
  nand GNAME6293(G6293,G1240,G21560);
  nand GNAME6294(G6294,G1661,G7714);
  nand GNAME6295(G6295,G6275,G1662);
  nand GNAME6296(G6296,G6292,G1687);
  nand GNAME6297(G6297,G6258,G1260);
  nand GNAME6298(G6298,G21556,G1691);
  nand GNAME6299(G6299,G21548,G1693);
  nand GNAME6300(G6300,G21540,G1695);
  nand GNAME6301(G6301,G21532,G1696);
  nand GNAME6302(G6302,G21524,G1698);
  nand GNAME6303(G6303,G21516,G1700);
  nand GNAME6304(G6304,G21508,G1701);
  nand GNAME6305(G6305,G21500,G1702);
  nand GNAME6306(G6306,G21492,G1704);
  nand GNAME6307(G6307,G21484,G1705);
  nand GNAME6308(G6308,G21476,G1707);
  nand GNAME6309(G6309,G21468,G1708);
  nand GNAME6310(G6310,G21460,G1709);
  nand GNAME6311(G6311,G21452,G1710);
  nand GNAME6312(G6312,G21444,G1711);
  nand GNAME6313(G6313,G21436,G1712);
  nand GNAME6314(G6314,G2233,G2234,G2235,G2236);
  nand GNAME6315(G6315,G21436,G2286);
  nand GNAME6316(G6316,G21444,G2285);
  nand GNAME6317(G6317,G21452,G2284);
  nand GNAME6318(G6318,G21460,G2283);
  nand GNAME6319(G6319,G21468,G2282);
  nand GNAME6320(G6320,G21476,G2281);
  nand GNAME6321(G6321,G21484,G2280);
  nand GNAME6322(G6322,G21492,G2279);
  nand GNAME6323(G6323,G21500,G2276);
  nand GNAME6324(G6324,G21508,G2275);
  nand GNAME6325(G6325,G21516,G2274);
  nand GNAME6326(G6326,G21524,G2273);
  nand GNAME6327(G6327,G21532,G2272);
  nand GNAME6328(G6328,G21540,G2271);
  nand GNAME6329(G6329,G21548,G2270);
  nand GNAME6330(G6330,G21556,G2269);
  nand GNAME6331(G6331,G2225,G2226,G2227,G2228);
  nand GNAME6332(G6332,G21436,G1665);
  nand GNAME6333(G6333,G21444,G1667);
  nand GNAME6334(G6334,G21452,G1669);
  nand GNAME6335(G6335,G21460,G1670);
  nand GNAME6336(G6336,G21468,G1672);
  nand GNAME6337(G6337,G21476,G1674);
  nand GNAME6338(G6338,G21484,G1675);
  nand GNAME6339(G6339,G21492,G1676);
  nand GNAME6340(G6340,G21500,G1678);
  nand GNAME6341(G6341,G21508,G1679);
  nand GNAME6342(G6342,G21516,G1681);
  nand GNAME6343(G6343,G21524,G1682);
  nand GNAME6344(G6344,G21532,G1683);
  nand GNAME6345(G6345,G21540,G1684);
  nand GNAME6346(G6346,G21548,G1685);
  nand GNAME6347(G6347,G21556,G1686);
  nand GNAME6348(G6348,G2229,G2230,G2231,G2232);
  nand GNAME6349(G6349,G1240,G21561);
  nand GNAME6350(G6350,G1661,G7717);
  nand GNAME6351(G6351,G6331,G1662);
  nand GNAME6352(G6352,G6348,G1687);
  nand GNAME6353(G6353,G6314,G1260);
  nand GNAME6354(G6354,G21554,G1571);
  or GNAME6355(G6355,G1515,G2528,G1269);
  nand GNAME6356(G6356,G1243,G1253,G21428,G7294);
  nand GNAME6357(G6357,G21555,G1571);
  nand GNAME6358(G6358,G2511,G1253);
  nand GNAME6359(G6359,G1240,G2477);
  nand GNAME6360(G6360,G1282,G1511);
  nand GNAME6361(G6361,G1265,G1501);
  nand GNAME6362(G6362,G2239,G7279,G6360,G1520,G1716);
  nand GNAME6363(G6363,G6362,G21428);
  nand GNAME6364(G6364,G21556,G1571);
  nand GNAME6365(G6365,G1248,G1249);
  nand GNAME6366(G6366,G682,G1239);
  nand GNAME6367(G6367,G6366,G2600);
  nand GNAME6368(G6368,G1518,G1248,G1252);
  nand GNAME6369(G6369,G6367,G1501);
  nand GNAME6370(G6370,G6365,G1261);
  or GNAME6371(G6371,G2477,G1297);
  nand GNAME6372(G6372,G5209,G1509);
  nand GNAME6373(G6373,G2240,G6370,G6371,G6372,G1521);
  nand GNAME6374(G6374,G6373,G21428);
  or GNAME6375(G6375,G1269,G1717);
  or GNAME6376(G6376,G2511,G1718);
  nand GNAME6377(G6377,G2241,G1719,G6375,G2304);
  or GNAME6378(G6378,G1571,G1278);
  nand GNAME6379(G6379,G6378,G7468);
  nand GNAME6380(G6380,G4406,G21608);
  nand GNAME6381(G6381,G6377,G21576);
  nand GNAME6382(G6382,G21767,G2297);
  nand GNAME6383(G6383,G6378,G7469);
  nand GNAME6384(G6384,G4406,G21607);
  nand GNAME6385(G6385,G6377,G21575);
  nand GNAME6386(G6386,G21766,G2297);
  nand GNAME6387(G6387,G6378,G7445);
  nand GNAME6388(G6388,G4406,G21606);
  nand GNAME6389(G6389,G6377,G21574);
  nand GNAME6390(G6390,G21765,G2297);
  nand GNAME6391(G6391,G6378,G7444);
  nand GNAME6392(G6392,G4406,G21605);
  nand GNAME6393(G6393,G6377,G21573);
  nand GNAME6394(G6394,G21764,G2297);
  nand GNAME6395(G6395,G6378,G7470);
  nand GNAME6396(G6396,G4406,G21604);
  nand GNAME6397(G6397,G6377,G21572);
  nand GNAME6398(G6398,G21763,G2297);
  nand GNAME6399(G6399,G1557,G2303);
  nand GNAME6400(G6400,G6399,G21557);
  nand GNAME6401(G6401,G6378,G7471);
  nand GNAME6402(G6402,G4406,G21603);
  nand GNAME6403(G6403,G6377,G21571);
  nand GNAME6404(G6404,G21762,G2297);
  nand GNAME6405(G6405,G4406,G21630);
  nand GNAME6406(G6406,G6377,G21598);
  nand GNAME6407(G6407,G21789,G2297);
  nand GNAME6408(G6408,G1278,G7442);
  nand GNAME6409(G6409,G6378,G7441);
  nand GNAME6410(G6410,G4406,G21629);
  nand GNAME6411(G6411,G6377,G21597);
  nand GNAME6412(G6412,G21788,G2297);
  nand GNAME6413(G6413,G5492,G2300);
  nand GNAME6414(G6414,G2327,G2323,G2324);
  nand GNAME6415(G6415,G6414,G21428);
  or GNAME6416(G6416,G1248,G1718);
  or GNAME6417(G6417,G2545,G1720);
  nand GNAME6418(G6418,G2242,G1721,G6416,G6417);
  nand GNAME6419(G6419,G6418,G21558);
  nand GNAME6420(G6420,G6378,G7443);
  nand GNAME6421(G6421,G4406,G21602);
  nand GNAME6422(G6422,G6377,G21570);
  nand GNAME6423(G6423,G21761,G2297);
  nand GNAME6424(G6424,G6378,G7472);
  nand GNAME6425(G6425,G4406,G21628);
  nand GNAME6426(G6426,G6377,G21596);
  nand GNAME6427(G6427,G21787,G2297);
  nand GNAME6428(G6428,G5509,G2300);
  nand GNAME6429(G6429,G6378,G7473);
  nand GNAME6430(G6430,G4406,G21627);
  nand GNAME6431(G6431,G6377,G21595);
  nand GNAME6432(G6432,G21786,G2297);
  nand GNAME6433(G6433,G5526,G2300);
  nand GNAME6434(G6434,G6378,G7474);
  nand GNAME6435(G6435,G4406,G21626);
  nand GNAME6436(G6436,G6377,G21594);
  nand GNAME6437(G6437,G21785,G2297);
  nand GNAME6438(G6438,G5543,G2300);
  nand GNAME6439(G6439,G6378,G7475);
  nand GNAME6440(G6440,G4406,G21625);
  nand GNAME6441(G6441,G6377,G21593);
  nand GNAME6442(G6442,G21784,G2297);
  nand GNAME6443(G6443,G5560,G2300);
  nand GNAME6444(G6444,G6378,G7476);
  nand GNAME6445(G6445,G4406,G21624);
  nand GNAME6446(G6446,G6377,G21592);
  nand GNAME6447(G6447,G21783,G2297);
  nand GNAME6448(G6448,G5577,G2300);
  nand GNAME6449(G6449,G6378,G7477);
  nand GNAME6450(G6450,G4406,G21623);
  nand GNAME6451(G6451,G6377,G21591);
  nand GNAME6452(G6452,G21782,G2297);
  nand GNAME6453(G6453,G5594,G2300);
  nand GNAME6454(G6454,G6378,G7478);
  nand GNAME6455(G6455,G4406,G21622);
  nand GNAME6456(G6456,G6377,G21590);
  nand GNAME6457(G6457,G21781,G2297);
  nand GNAME6458(G6458,G5611,G2300);
  nand GNAME6459(G6459,G6378,G7479);
  nand GNAME6460(G6460,G4406,G21621);
  nand GNAME6461(G6461,G6377,G21589);
  nand GNAME6462(G6462,G21780,G2297);
  nand GNAME6463(G6463,G6378,G7480);
  nand GNAME6464(G6464,G4406,G21620);
  nand GNAME6465(G6465,G6377,G21588);
  nand GNAME6466(G6466,G21779,G2297);
  nand GNAME6467(G6467,G6378,G7481);
  nand GNAME6468(G6468,G4406,G21619);
  nand GNAME6469(G6469,G6377,G21587);
  nand GNAME6470(G6470,G21778,G2297);
  nand GNAME6471(G6471,G6418,G21559);
  nand GNAME6472(G6472,G6378,G7440);
  nand GNAME6473(G6473,G4406,G21601);
  nand GNAME6474(G6474,G6377,G21569);
  nand GNAME6475(G6475,G21760,G2297);
  nand GNAME6476(G6476,G6378,G7483);
  nand GNAME6477(G6477,G4406,G21618);
  nand GNAME6478(G6478,G6377,G21586);
  nand GNAME6479(G6479,G21777,G2297);
  nand GNAME6480(G6480,G6378,G7484);
  nand GNAME6481(G6481,G4406,G21617);
  nand GNAME6482(G6482,G6377,G21585);
  nand GNAME6483(G6483,G21776,G2297);
  nand GNAME6484(G6484,G6378,G7485);
  nand GNAME6485(G6485,G4406,G21616);
  nand GNAME6486(G6486,G6377,G21584);
  nand GNAME6487(G6487,G21775,G2297);
  nand GNAME6488(G6488,G6378,G7486);
  nand GNAME6489(G6489,G4406,G21615);
  nand GNAME6490(G6490,G6377,G21583);
  nand GNAME6491(G6491,G21774,G2297);
  nand GNAME6492(G6492,G6378,G7487);
  nand GNAME6493(G6493,G4406,G21614);
  nand GNAME6494(G6494,G6377,G21582);
  nand GNAME6495(G6495,G21773,G2297);
  nand GNAME6496(G6496,G6378,G7439);
  nand GNAME6497(G6497,G4406,G21613);
  nand GNAME6498(G6498,G6377,G21581);
  nand GNAME6499(G6499,G21772,G2297);
  nand GNAME6500(G6500,G6378,G7488);
  nand GNAME6501(G6501,G4406,G21612);
  nand GNAME6502(G6502,G6377,G21580);
  nand GNAME6503(G6503,G21771,G2297);
  nand GNAME6504(G6504,G6378,G7489);
  nand GNAME6505(G6505,G4406,G21611);
  nand GNAME6506(G6506,G6377,G21579);
  nand GNAME6507(G6507,G21770,G2297);
  nand GNAME6508(G6508,G6378,G7438);
  nand GNAME6509(G6509,G4406,G21610);
  nand GNAME6510(G6510,G6377,G21578);
  nand GNAME6511(G6511,G21769,G2297);
  nand GNAME6512(G6512,G6378,G7437);
  nand GNAME6513(G6513,G4406,G21609);
  nand GNAME6514(G6514,G6377,G21577);
  nand GNAME6515(G6515,G21768,G2297);
  nand GNAME6516(G6516,G6418,G21560);
  nand GNAME6517(G6517,G6378,G7482);
  nand GNAME6518(G6518,G4406,G21600);
  nand GNAME6519(G6519,G6377,G21568);
  nand GNAME6520(G6520,G21759,G2297);
  nand GNAME6521(G6521,G6418,G21561);
  nand GNAME6522(G6522,G6378,G7467);
  nand GNAME6523(G6523,G4406,G21599);
  nand GNAME6524(G6524,G6377,G21567);
  nand GNAME6525(G6525,G21758,G2297);
  nand GNAME6526(G6526,G7284,G2579);
  nand GNAME6527(G6527,G2596,G1265);
  nand GNAME6528(G6528,G1238,G1501);
  nand GNAME6529(G6529,G2243,G7281,G7282,G6752,G1716);
  nand GNAME6530(G6530,G6529,G21428);
  nand GNAME6531(G6531,G2301,G1720,G1718,G1721);
  nand GNAME6532(G6532,G2299,G1551);
  nand GNAME6533(G6533,G6532,G21735);
  nand GNAME6534(G6534,G6531,G21576);
  nand GNAME6535(G6535,G21703,G2302);
  nand GNAME6536(G6536,G8754,G1571);
  nand GNAME6537(G6537,G1278,G21608);
  nand GNAME6538(G6538,G6532,G21734);
  nand GNAME6539(G6539,G6531,G21575);
  nand GNAME6540(G6540,G21702,G2302);
  nand GNAME6541(G6541,G8755,G1571);
  nand GNAME6542(G6542,G1278,G21607);
  nand GNAME6543(G6543,G6532,G21733);
  nand GNAME6544(G6544,G6531,G21574);
  nand GNAME6545(G6545,G21701,G2302);
  nand GNAME6546(G6546,G8756,G1571);
  nand GNAME6547(G6547,G1278,G21606);
  nand GNAME6548(G6548,G6532,G21732);
  nand GNAME6549(G6549,G6531,G21573);
  nand GNAME6550(G6550,G21700,G2302);
  nand GNAME6551(G6551,G8757,G1571);
  nand GNAME6552(G6552,G1278,G21605);
  nand GNAME6553(G6553,G6532,G21731);
  nand GNAME6554(G6554,G6531,G21572);
  nand GNAME6555(G6555,G21699,G2302);
  nand GNAME6556(G6556,G8758,G1571);
  nand GNAME6557(G6557,G1278,G21604);
  nand GNAME6558(G6558,G6532,G21730);
  nand GNAME6559(G6559,G6531,G21571);
  nand GNAME6560(G6560,G21698,G2302);
  nand GNAME6561(G6561,G8759,G1571);
  nand GNAME6562(G6562,G1278,G21603);
  nand GNAME6563(G6563,G6532,G21757);
  nand GNAME6564(G6564,G6531,G21598);
  nand GNAME6565(G6565,G21725,G2302);
  nand GNAME6566(G6566,G1278,G21630);
  nand GNAME6567(G6567,G6532,G21756);
  nand GNAME6568(G6568,G6531,G21597);
  nand GNAME6569(G6569,G21724,G2302);
  nand GNAME6570(G6570,G8760,G1571);
  nand GNAME6571(G6571,G1278,G21629);
  nand GNAME6572(G6572,G1719,G1713,G1714);
  nand GNAME6573(G6573,G6572,G21558);
  nand GNAME6574(G6574,G6532,G21729);
  nand GNAME6575(G6575,G6531,G21570);
  nand GNAME6576(G6576,G1281,G21563);
  nand GNAME6577(G6577,G21697,G2302);
  nand GNAME6578(G6578,G8782,G1571);
  nand GNAME6579(G6579,G1278,G21602);
  nand GNAME6580(G6580,G1729,G1277);
  nand GNAME6581(G6581,G1292,G6804);
  nand GNAME6582(G6582,G6532,G21755);
  nand GNAME6583(G6583,G6531,G21596);
  nand GNAME6584(G6584,G21723,G2302);
  nand GNAME6585(G6585,G8707,G1571);
  nand GNAME6586(G6586,G1278,G21628);
  nand GNAME6587(G6587,G6532,G21754);
  nand GNAME6588(G6588,G6531,G21595);
  nand GNAME6589(G6589,G21722,G2302);
  nand GNAME6590(G6590,G8706,G1571);
  nand GNAME6591(G6591,G1278,G21627);
  nand GNAME6592(G6592,G6532,G21753);
  nand GNAME6593(G6593,G6531,G21594);
  nand GNAME6594(G6594,G21721,G2302);
  nand GNAME6595(G6595,G8761,G1571);
  nand GNAME6596(G6596,G1278,G21626);
  nand GNAME6597(G6597,G6532,G21752);
  nand GNAME6598(G6598,G6531,G21593);
  nand GNAME6599(G6599,G21720,G2302);
  nand GNAME6600(G6600,G8705,G1571);
  nand GNAME6601(G6601,G1278,G21625);
  nand GNAME6602(G6602,G6532,G21751);
  nand GNAME6603(G6603,G6531,G21592);
  nand GNAME6604(G6604,G21719,G2302);
  nand GNAME6605(G6605,G8704,G1571);
  nand GNAME6606(G6606,G1278,G21624);
  nand GNAME6607(G6607,G6532,G21750);
  nand GNAME6608(G6608,G6531,G21591);
  nand GNAME6609(G6609,G21718,G2302);
  nand GNAME6610(G6610,G8785,G1571);
  nand GNAME6611(G6611,G1278,G21623);
  nand GNAME6612(G6612,G6532,G21749);
  nand GNAME6613(G6613,G6531,G21590);
  nand GNAME6614(G6614,G21717,G2302);
  nand GNAME6615(G6615,G8771,G1571);
  nand GNAME6616(G6616,G1278,G21622);
  nand GNAME6617(G6617,G6532,G21748);
  nand GNAME6618(G6618,G6531,G21589);
  nand GNAME6619(G6619,G21716,G2302);
  nand GNAME6620(G6620,G8772,G1571);
  nand GNAME6621(G6621,G1278,G21621);
  nand GNAME6622(G6622,G6532,G21747);
  nand GNAME6623(G6623,G6531,G21588);
  nand GNAME6624(G6624,G21715,G2302);
  nand GNAME6625(G6625,G8773,G1571);
  nand GNAME6626(G6626,G1278,G21620);
  nand GNAME6627(G6627,G6532,G21746);
  nand GNAME6628(G6628,G6531,G21587);
  nand GNAME6629(G6629,G21714,G2302);
  nand GNAME6630(G6630,G8774,G1571);
  nand GNAME6631(G6631,G1278,G21619);
  nand GNAME6632(G6632,G6572,G21559);
  nand GNAME6633(G6633,G6532,G21728);
  nand GNAME6634(G6634,G6531,G21569);
  nand GNAME6635(G6635,G1281,G21564);
  nand GNAME6636(G6636,G21696,G2302);
  nand GNAME6637(G6637,G8708,G1571);
  nand GNAME6638(G6638,G1278,G21601);
  nand GNAME6639(G6639,G1277,G1739);
  nand GNAME6640(G6640,G1292,G2259);
  nand GNAME6641(G6641,G6532,G21745);
  nand GNAME6642(G6642,G6531,G21586);
  nand GNAME6643(G6643,G21713,G2302);
  nand GNAME6644(G6644,G8775,G1571);
  nand GNAME6645(G6645,G1278,G21618);
  nand GNAME6646(G6646,G6532,G21744);
  nand GNAME6647(G6647,G6531,G21585);
  nand GNAME6648(G6648,G21712,G2302);
  nand GNAME6649(G6649,G8776,G1571);
  nand GNAME6650(G6650,G1278,G21617);
  nand GNAME6651(G6651,G6532,G21743);
  nand GNAME6652(G6652,G6531,G21584);
  nand GNAME6653(G6653,G21711,G2302);
  nand GNAME6654(G6654,G8777,G1571);
  nand GNAME6655(G6655,G1278,G21616);
  nand GNAME6656(G6656,G6532,G21742);
  nand GNAME6657(G6657,G6531,G21583);
  nand GNAME6658(G6658,G21710,G2302);
  nand GNAME6659(G6659,G8763,G1571);
  nand GNAME6660(G6660,G1278,G21615);
  nand GNAME6661(G6661,G6532,G21741);
  nand GNAME6662(G6662,G6531,G21582);
  nand GNAME6663(G6663,G21709,G2302);
  nand GNAME6664(G6664,G8764,G1571);
  nand GNAME6665(G6665,G1278,G21614);
  nand GNAME6666(G6666,G6532,G21740);
  nand GNAME6667(G6667,G6531,G21581);
  nand GNAME6668(G6668,G21708,G2302);
  nand GNAME6669(G6669,G8765,G1571);
  nand GNAME6670(G6670,G1278,G21613);
  nand GNAME6671(G6671,G6532,G21739);
  nand GNAME6672(G6672,G6531,G21580);
  nand GNAME6673(G6673,G21707,G2302);
  nand GNAME6674(G6674,G8766,G1571);
  nand GNAME6675(G6675,G1278,G21612);
  nand GNAME6676(G6676,G6532,G21738);
  nand GNAME6677(G6677,G6531,G21579);
  nand GNAME6678(G6678,G21706,G2302);
  nand GNAME6679(G6679,G8767,G1571);
  nand GNAME6680(G6680,G1278,G21611);
  nand GNAME6681(G6681,G6532,G21737);
  nand GNAME6682(G6682,G6531,G21578);
  nand GNAME6683(G6683,G21705,G2302);
  nand GNAME6684(G6684,G8768,G1571);
  nand GNAME6685(G6685,G1278,G21610);
  nand GNAME6686(G6686,G6532,G21736);
  nand GNAME6687(G6687,G6531,G21577);
  nand GNAME6688(G6688,G21704,G2302);
  nand GNAME6689(G6689,G8769,G1571);
  nand GNAME6690(G6690,G1278,G21609);
  nand GNAME6691(G6691,G6572,G21560);
  nand GNAME6692(G6692,G6532,G21727);
  nand GNAME6693(G6693,G6531,G21568);
  nand GNAME6694(G6694,G1281,G21565);
  nand GNAME6695(G6695,G21695,G2302);
  nand GNAME6696(G6696,G8762,G1571);
  nand GNAME6697(G6697,G1278,G21600);
  nand GNAME6698(G6698,G1728,G1277);
  nand GNAME6699(G6699,G1727,G1292);
  nand GNAME6700(G6700,G6572,G21561);
  nand GNAME6701(G6701,G6532,G21726);
  nand GNAME6702(G6702,G6531,G21567);
  nand GNAME6703(G6703,G1281,G21566);
  nand GNAME6704(G6704,G21694,G2302);
  nand GNAME6705(G6705,G8709,G1571);
  nand GNAME6706(G6706,G1278,G21599);
  nand GNAME6707(G6707,G1277,G2277);
  nand GNAME6708(G6708,G1292,G2258);
  nand GNAME6709(G6709,G6107,G2296);
  or GNAME6710(G6710,G1208,G7289);
  nand GNAME6711(G6711,G6163,G2296);
  nand GNAME6712(G6712,G21425,G21558);
  nand GNAME6713(G6713,G1280,G1242,G2528);
  nand GNAME6714(G6714,G6219,G2296);
  nand GNAME6715(G6715,G21425,G21559);
  nand GNAME6716(G6716,G1242,G7283,G7284);
  nand GNAME6717(G6717,G6275,G2296);
  nand GNAME6718(G6718,G1242,G2528);
  nand GNAME6719(G6719,G6718,G2329);
  nand GNAME6720(G6720,G6331,G2296);
  nand GNAME6721(G6721,G1238,G1242,G1249);
  nand GNAME6722(G6722,G6721,G1280);
  nand GNAME6723(G6723,G6722,G2295);
  nand GNAME6724(G6724,G6723,G8132);
  nand GNAME6725(G6725,G6723,G8149);
  nand GNAME6726(G6726,G21427,G558);
  nand GNAME6727(G6727,G6723,G8151);
  nand GNAME6728(G6728,G21427,G8702);
  nand GNAME6729(G6729,G6723,G8153);
  nand GNAME6730(G6730,G21427,G8703);
  nand GNAME6731(G6731,G6723,G8143);
  nand GNAME6732(G6732,G21427,G8700);
  nand GNAME6733(G6733,G6723,G8133);
  nand GNAME6734(G6734,G21427,G8701);
  nand GNAME6735(G6735,G1511,G1242,G1249);
  nand GNAME6736(G6736,G1208,G6735);
  nand GNAME6737(G6737,G4997,G1578);
  nand GNAME6738(G6738,G1300,G1579);
  nand GNAME6739(G6739,G1760,G1579);
  nand GNAME6740(G6740,G6738,G2334,G6737);
  nand GNAME6741(G6741,G2331,G6739);
  or GNAME6742(G6742,G2337,G1584);
  nand GNAME6743(G6743,G21391,G2315,G2316);
  nand GNAME6744(G6744,G21392,G2314,G2316);
  nand GNAME6745(G6745,G1197,G2316);
  nand GNAME6746(G6746,G1240,G2599);
  or GNAME6747(G6747,G8101,G1190);
  or GNAME6748(G6748,G2611,G1257);
  nor GNAME6749(G6749,G1208,G1271);
  nand GNAME6750(G6750,G1252,G2562);
  nand GNAME6751(G6751,G21393,G21758);
  nand GNAME6752(G6752,G2528,G1516);
  nand GNAME6753(G6753,G2313,G21356);
  nand GNAME6754(G6754,G1195,G21790);
  nand GNAME6755(G6755,G2313,G21357);
  nand GNAME6756(G6756,G1195,G21791);
  nand GNAME6757(G6757,G2313,G21358);
  nand GNAME6758(G6758,G1195,G21792);
  nand GNAME6759(G6759,G2313,G21359);
  nand GNAME6760(G6760,G1195,G21793);
  or GNAME6761(G6761,G33,G21392);
  nand GNAME6762(G6762,G21392,G788,G1205);
  nand GNAME6763(G6763,G1204,G21390);
  nand GNAME6764(G6764,G21392,G2453,G21798);
  nand GNAME6765(G6765,G6763,G6764);
  nand GNAME6766(G6766,G2450,G21391);
  nand GNAME6767(G6767,G1194,G6765);
  and GNAME6768(G6768,G2454,G21392);
  and GNAME6769(G6769,G1204,G2456);
  or GNAME6770(G6770,G21391,G21392);
  nand GNAME6771(G6771,G1201,G21392);
  not GNAME6772(G6772,G1736);
  nand GNAME6773(G6773,G21393,G6772);
  or GNAME6774(G6774,G6772,G34,G1589);
  nand GNAME6775(G6775,G2457,G1736);
  nand GNAME6776(G6776,G21394,G6772);
  or GNAME6777(G6777,G21428,G35);
  nand GNAME6778(G6778,G2613,G21428);
  or GNAME6779(G6779,G1269,G1271);
  nand GNAME6780(G6780,G1271,G2627);
  nand GNAME6781(G6781,G1272,G1292);
  nand GNAME6782(G6782,G21427,G1269,G1209);
  or GNAME6783(G6783,G21426,G21566);
  nand GNAME6784(G6784,G21566,G1292);
  nand GNAME6785(G6785,G1300,G21567);
  nand GNAME6786(G6786,G1760,G21567);
  nand GNAME6787(G6787,G6785,G6786);
  or GNAME6788(G6788,G21568,G1760);
  or GNAME6789(G6789,G1300,G7297);
  nand GNAME6790(G6790,G1305,G2634);
  nand GNAME6791(G6791,G1304,G2646);
  nand GNAME6792(G6792,G1306,G1802);
  or GNAME6793(G6793,G1306,G1802);
  not GNAME6794(G6794,G1727);
  nand GNAME6795(G6795,G2683,G2677);
  nand GNAME6796(G6796,G1311,G2681,G2682);
  nand GNAME6797(G6797,G1307,G2656);
  nand GNAME6798(G6798,G1298,G2669);
  nand GNAME6799(G6799,G2673,G1803);
  or GNAME6800(G6800,G2673,G1803);
  not GNAME6801(G6801,G1728);
  nand GNAME6802(G6802,G2249,G2248);
  or GNAME6803(G6803,G2248,G2249);
  not GNAME6804(G6804,G1726);
  nand GNAME6805(G6805,G2251,G2250);
  or GNAME6806(G6806,G2250,G2251);
  not GNAME6807(G6807,G1729);
  nand GNAME6808(G6808,G2294,G21429);
  nand GNAME6809(G6809,G1294,G25);
  nand GNAME6810(G6810,G6808,G6809);
  nand GNAME6811(G6811,G2294,G21430);
  nand GNAME6812(G6812,G1294,G26);
  nand GNAME6813(G6813,G6811,G6812);
  nand GNAME6814(G6814,G2294,G21431);
  nand GNAME6815(G6815,G1294,G27);
  nand GNAME6816(G6816,G6814,G6815);
  nand GNAME6817(G6817,G2294,G21432);
  nand GNAME6818(G6818,G1294,G28);
  nand GNAME6819(G6819,G6817,G6818);
  nand GNAME6820(G6820,G2294,G21433);
  nand GNAME6821(G6821,G1294,G29);
  nand GNAME6822(G6822,G6820,G6821);
  nand GNAME6823(G6823,G2294,G21434);
  nand GNAME6824(G6824,G1294,G30);
  nand GNAME6825(G6825,G6823,G6824);
  nand GNAME6826(G6826,G2294,G21435);
  nand GNAME6827(G6827,G1294,G31);
  nand GNAME6828(G6828,G6826,G6827);
  nand GNAME6829(G6829,G2294,G21436);
  nand GNAME6830(G6830,G1294,G32);
  nand GNAME6831(G6831,G6829,G6830);
  nand GNAME6832(G6832,G1353,G21437);
  nand GNAME6833(G6833,G25,G2293);
  nand GNAME6834(G6834,G6832,G6833);
  nand GNAME6835(G6835,G1353,G21438);
  nand GNAME6836(G6836,G26,G2293);
  nand GNAME6837(G6837,G6835,G6836);
  nand GNAME6838(G6838,G1353,G21439);
  nand GNAME6839(G6839,G27,G2293);
  nand GNAME6840(G6840,G6838,G6839);
  nand GNAME6841(G6841,G1353,G21440);
  nand GNAME6842(G6842,G28,G2293);
  nand GNAME6843(G6843,G6841,G6842);
  nand GNAME6844(G6844,G1353,G21441);
  nand GNAME6845(G6845,G29,G2293);
  nand GNAME6846(G6846,G6844,G6845);
  nand GNAME6847(G6847,G1353,G21442);
  nand GNAME6848(G6848,G30,G2293);
  nand GNAME6849(G6849,G6847,G6848);
  nand GNAME6850(G6850,G1353,G21443);
  nand GNAME6851(G6851,G31,G2293);
  nand GNAME6852(G6852,G6850,G6851);
  nand GNAME6853(G6853,G1353,G21444);
  nand GNAME6854(G6854,G32,G2293);
  nand GNAME6855(G6855,G6853,G6854);
  nand GNAME6856(G6856,G1367,G21445);
  nand GNAME6857(G6857,G25,G2292);
  nand GNAME6858(G6858,G6856,G6857);
  nand GNAME6859(G6859,G1367,G21446);
  nand GNAME6860(G6860,G26,G2292);
  nand GNAME6861(G6861,G6859,G6860);
  nand GNAME6862(G6862,G1367,G21447);
  nand GNAME6863(G6863,G27,G2292);
  nand GNAME6864(G6864,G6862,G6863);
  nand GNAME6865(G6865,G1367,G21448);
  nand GNAME6866(G6866,G28,G2292);
  nand GNAME6867(G6867,G6865,G6866);
  nand GNAME6868(G6868,G1367,G21449);
  nand GNAME6869(G6869,G29,G2292);
  nand GNAME6870(G6870,G6868,G6869);
  nand GNAME6871(G6871,G1367,G21450);
  nand GNAME6872(G6872,G30,G2292);
  nand GNAME6873(G6873,G6871,G6872);
  nand GNAME6874(G6874,G1367,G21451);
  nand GNAME6875(G6875,G31,G2292);
  nand GNAME6876(G6876,G6874,G6875);
  nand GNAME6877(G6877,G1367,G21452);
  nand GNAME6878(G6878,G32,G2292);
  nand GNAME6879(G6879,G6877,G6878);
  nand GNAME6880(G6880,G1379,G21453);
  nand GNAME6881(G6881,G25,G2291);
  nand GNAME6882(G6882,G6880,G6881);
  nand GNAME6883(G6883,G1379,G21454);
  nand GNAME6884(G6884,G26,G2291);
  nand GNAME6885(G6885,G6883,G6884);
  nand GNAME6886(G6886,G1379,G21455);
  nand GNAME6887(G6887,G27,G2291);
  nand GNAME6888(G6888,G6886,G6887);
  nand GNAME6889(G6889,G1379,G21456);
  nand GNAME6890(G6890,G28,G2291);
  nand GNAME6891(G6891,G6889,G6890);
  nand GNAME6892(G6892,G1379,G21457);
  nand GNAME6893(G6893,G29,G2291);
  nand GNAME6894(G6894,G6892,G6893);
  nand GNAME6895(G6895,G1379,G21458);
  nand GNAME6896(G6896,G30,G2291);
  nand GNAME6897(G6897,G6895,G6896);
  nand GNAME6898(G6898,G1379,G21459);
  nand GNAME6899(G6899,G31,G2291);
  nand GNAME6900(G6900,G6898,G6899);
  nand GNAME6901(G6901,G1379,G21460);
  nand GNAME6902(G6902,G32,G2291);
  nand GNAME6903(G6903,G6901,G6902);
  nand GNAME6904(G6904,G1391,G21461);
  nand GNAME6905(G6905,G25,G2290);
  nand GNAME6906(G6906,G6904,G6905);
  nand GNAME6907(G6907,G1391,G21462);
  nand GNAME6908(G6908,G26,G2290);
  nand GNAME6909(G6909,G6907,G6908);
  nand GNAME6910(G6910,G1391,G21463);
  nand GNAME6911(G6911,G27,G2290);
  nand GNAME6912(G6912,G6910,G6911);
  nand GNAME6913(G6913,G1391,G21464);
  nand GNAME6914(G6914,G28,G2290);
  nand GNAME6915(G6915,G6913,G6914);
  nand GNAME6916(G6916,G1391,G21465);
  nand GNAME6917(G6917,G29,G2290);
  nand GNAME6918(G6918,G6916,G6917);
  nand GNAME6919(G6919,G1391,G21466);
  nand GNAME6920(G6920,G30,G2290);
  nand GNAME6921(G6921,G6919,G6920);
  nand GNAME6922(G6922,G1391,G21467);
  nand GNAME6923(G6923,G31,G2290);
  nand GNAME6924(G6924,G6922,G6923);
  nand GNAME6925(G6925,G1391,G21468);
  nand GNAME6926(G6926,G32,G2290);
  nand GNAME6927(G6927,G6925,G6926);
  nand GNAME6928(G6928,G1402,G21469);
  nand GNAME6929(G6929,G25,G2289);
  nand GNAME6930(G6930,G6928,G6929);
  nand GNAME6931(G6931,G1402,G21470);
  nand GNAME6932(G6932,G26,G2289);
  nand GNAME6933(G6933,G6931,G6932);
  nand GNAME6934(G6934,G1402,G21471);
  nand GNAME6935(G6935,G27,G2289);
  nand GNAME6936(G6936,G6934,G6935);
  nand GNAME6937(G6937,G1402,G21472);
  nand GNAME6938(G6938,G28,G2289);
  nand GNAME6939(G6939,G6937,G6938);
  nand GNAME6940(G6940,G1402,G21473);
  nand GNAME6941(G6941,G29,G2289);
  nand GNAME6942(G6942,G6940,G6941);
  nand GNAME6943(G6943,G1402,G21474);
  nand GNAME6944(G6944,G30,G2289);
  nand GNAME6945(G6945,G6943,G6944);
  nand GNAME6946(G6946,G1402,G21475);
  nand GNAME6947(G6947,G31,G2289);
  nand GNAME6948(G6948,G6946,G6947);
  nand GNAME6949(G6949,G1402,G21476);
  nand GNAME6950(G6950,G32,G2289);
  nand GNAME6951(G6951,G6949,G6950);
  nand GNAME6952(G6952,G1413,G21477);
  nand GNAME6953(G6953,G25,G2288);
  nand GNAME6954(G6954,G6952,G6953);
  nand GNAME6955(G6955,G1413,G21478);
  nand GNAME6956(G6956,G26,G2288);
  nand GNAME6957(G6957,G6955,G6956);
  nand GNAME6958(G6958,G1413,G21479);
  nand GNAME6959(G6959,G27,G2288);
  nand GNAME6960(G6960,G6958,G6959);
  nand GNAME6961(G6961,G1413,G21480);
  nand GNAME6962(G6962,G28,G2288);
  nand GNAME6963(G6963,G6961,G6962);
  nand GNAME6964(G6964,G1413,G21481);
  nand GNAME6965(G6965,G29,G2288);
  nand GNAME6966(G6966,G6964,G6965);
  nand GNAME6967(G6967,G1413,G21482);
  nand GNAME6968(G6968,G30,G2288);
  nand GNAME6969(G6969,G6967,G6968);
  nand GNAME6970(G6970,G1413,G21483);
  nand GNAME6971(G6971,G31,G2288);
  nand GNAME6972(G6972,G6970,G6971);
  nand GNAME6973(G6973,G1413,G21484);
  nand GNAME6974(G6974,G32,G2288);
  nand GNAME6975(G6975,G6973,G6974);
  nand GNAME6976(G6976,G1423,G21485);
  nand GNAME6977(G6977,G25,G2287);
  nand GNAME6978(G6978,G6976,G6977);
  nand GNAME6979(G6979,G1423,G21486);
  nand GNAME6980(G6980,G26,G2287);
  nand GNAME6981(G6981,G6979,G6980);
  nand GNAME6982(G6982,G1423,G21487);
  nand GNAME6983(G6983,G27,G2287);
  nand GNAME6984(G6984,G6982,G6983);
  nand GNAME6985(G6985,G1423,G21488);
  nand GNAME6986(G6986,G28,G2287);
  nand GNAME6987(G6987,G6985,G6986);
  nand GNAME6988(G6988,G1423,G21489);
  nand GNAME6989(G6989,G29,G2287);
  nand GNAME6990(G6990,G6988,G6989);
  nand GNAME6991(G6991,G1423,G21490);
  nand GNAME6992(G6992,G30,G2287);
  nand GNAME6993(G6993,G6991,G6992);
  nand GNAME6994(G6994,G1423,G21491);
  nand GNAME6995(G6995,G31,G2287);
  nand GNAME6996(G6996,G6994,G6995);
  nand GNAME6997(G6997,G1423,G21492);
  nand GNAME6998(G6998,G32,G2287);
  nand GNAME6999(G6999,G6997,G6998);
  nand GNAME7000(G7000,G2268,G21493);
  nand GNAME7001(G7001,G25,G1435);
  nand GNAME7002(G7002,G7000,G7001);
  nand GNAME7003(G7003,G2268,G21494);
  nand GNAME7004(G7004,G26,G1435);
  nand GNAME7005(G7005,G7003,G7004);
  nand GNAME7006(G7006,G2268,G21495);
  nand GNAME7007(G7007,G27,G1435);
  nand GNAME7008(G7008,G7006,G7007);
  nand GNAME7009(G7009,G2268,G21496);
  nand GNAME7010(G7010,G28,G1435);
  nand GNAME7011(G7011,G7009,G7010);
  nand GNAME7012(G7012,G2268,G21497);
  nand GNAME7013(G7013,G29,G1435);
  nand GNAME7014(G7014,G7012,G7013);
  nand GNAME7015(G7015,G2268,G21498);
  nand GNAME7016(G7016,G30,G1435);
  nand GNAME7017(G7017,G7015,G7016);
  nand GNAME7018(G7018,G2268,G21499);
  nand GNAME7019(G7019,G31,G1435);
  nand GNAME7020(G7020,G7018,G7019);
  nand GNAME7021(G7021,G2268,G21500);
  nand GNAME7022(G7022,G32,G1435);
  nand GNAME7023(G7023,G7021,G7022);
  nand GNAME7024(G7024,G1443,G21501);
  nand GNAME7025(G7025,G25,G2267);
  nand GNAME7026(G7026,G7024,G7025);
  nand GNAME7027(G7027,G1443,G21502);
  nand GNAME7028(G7028,G26,G2267);
  nand GNAME7029(G7029,G7027,G7028);
  nand GNAME7030(G7030,G1443,G21503);
  nand GNAME7031(G7031,G27,G2267);
  nand GNAME7032(G7032,G7030,G7031);
  nand GNAME7033(G7033,G1443,G21504);
  nand GNAME7034(G7034,G28,G2267);
  nand GNAME7035(G7035,G7033,G7034);
  nand GNAME7036(G7036,G1443,G21505);
  nand GNAME7037(G7037,G29,G2267);
  nand GNAME7038(G7038,G7036,G7037);
  nand GNAME7039(G7039,G1443,G21506);
  nand GNAME7040(G7040,G30,G2267);
  nand GNAME7041(G7041,G7039,G7040);
  nand GNAME7042(G7042,G1443,G21507);
  nand GNAME7043(G7043,G31,G2267);
  nand GNAME7044(G7044,G7042,G7043);
  nand GNAME7045(G7045,G1443,G21508);
  nand GNAME7046(G7046,G32,G2267);
  nand GNAME7047(G7047,G7045,G7046);
  nand GNAME7048(G7048,G1452,G21509);
  nand GNAME7049(G7049,G25,G2266);
  nand GNAME7050(G7050,G7048,G7049);
  nand GNAME7051(G7051,G1452,G21510);
  nand GNAME7052(G7052,G26,G2266);
  nand GNAME7053(G7053,G7051,G7052);
  nand GNAME7054(G7054,G1452,G21511);
  nand GNAME7055(G7055,G27,G2266);
  nand GNAME7056(G7056,G7054,G7055);
  nand GNAME7057(G7057,G1452,G21512);
  nand GNAME7058(G7058,G28,G2266);
  nand GNAME7059(G7059,G7057,G7058);
  nand GNAME7060(G7060,G1452,G21513);
  nand GNAME7061(G7061,G29,G2266);
  nand GNAME7062(G7062,G7060,G7061);
  nand GNAME7063(G7063,G1452,G21514);
  nand GNAME7064(G7064,G30,G2266);
  nand GNAME7065(G7065,G7063,G7064);
  nand GNAME7066(G7066,G1452,G21515);
  nand GNAME7067(G7067,G31,G2266);
  nand GNAME7068(G7068,G7066,G7067);
  nand GNAME7069(G7069,G1452,G21516);
  nand GNAME7070(G7070,G32,G2266);
  nand GNAME7071(G7071,G7069,G7070);
  nand GNAME7072(G7072,G1460,G21517);
  nand GNAME7073(G7073,G25,G2265);
  nand GNAME7074(G7074,G7072,G7073);
  nand GNAME7075(G7075,G1460,G21518);
  nand GNAME7076(G7076,G26,G2265);
  nand GNAME7077(G7077,G7075,G7076);
  nand GNAME7078(G7078,G1460,G21519);
  nand GNAME7079(G7079,G27,G2265);
  nand GNAME7080(G7080,G7078,G7079);
  nand GNAME7081(G7081,G1460,G21520);
  nand GNAME7082(G7082,G28,G2265);
  nand GNAME7083(G7083,G7081,G7082);
  nand GNAME7084(G7084,G1460,G21521);
  nand GNAME7085(G7085,G29,G2265);
  nand GNAME7086(G7086,G7084,G7085);
  nand GNAME7087(G7087,G1460,G21522);
  nand GNAME7088(G7088,G30,G2265);
  nand GNAME7089(G7089,G7087,G7088);
  nand GNAME7090(G7090,G1460,G21523);
  nand GNAME7091(G7091,G31,G2265);
  nand GNAME7092(G7092,G7090,G7091);
  nand GNAME7093(G7093,G1460,G21524);
  nand GNAME7094(G7094,G32,G2265);
  nand GNAME7095(G7095,G7093,G7094);
  nand GNAME7096(G7096,G1469,G21525);
  nand GNAME7097(G7097,G25,G2264);
  nand GNAME7098(G7098,G7096,G7097);
  nand GNAME7099(G7099,G1469,G21526);
  nand GNAME7100(G7100,G26,G2264);
  nand GNAME7101(G7101,G7099,G7100);
  nand GNAME7102(G7102,G1469,G21527);
  nand GNAME7103(G7103,G27,G2264);
  nand GNAME7104(G7104,G7102,G7103);
  nand GNAME7105(G7105,G1469,G21528);
  nand GNAME7106(G7106,G28,G2264);
  nand GNAME7107(G7107,G7105,G7106);
  nand GNAME7108(G7108,G1469,G21529);
  nand GNAME7109(G7109,G29,G2264);
  nand GNAME7110(G7110,G7108,G7109);
  nand GNAME7111(G7111,G1469,G21530);
  nand GNAME7112(G7112,G30,G2264);
  nand GNAME7113(G7113,G7111,G7112);
  nand GNAME7114(G7114,G1469,G21531);
  nand GNAME7115(G7115,G31,G2264);
  nand GNAME7116(G7116,G7114,G7115);
  nand GNAME7117(G7117,G1469,G21532);
  nand GNAME7118(G7118,G32,G2264);
  nand GNAME7119(G7119,G7117,G7118);
  nand GNAME7120(G7120,G1477,G21533);
  nand GNAME7121(G7121,G25,G2263);
  nand GNAME7122(G7122,G7120,G7121);
  nand GNAME7123(G7123,G1477,G21534);
  nand GNAME7124(G7124,G26,G2263);
  nand GNAME7125(G7125,G7123,G7124);
  nand GNAME7126(G7126,G1477,G21535);
  nand GNAME7127(G7127,G27,G2263);
  nand GNAME7128(G7128,G7126,G7127);
  nand GNAME7129(G7129,G1477,G21536);
  nand GNAME7130(G7130,G28,G2263);
  nand GNAME7131(G7131,G7129,G7130);
  nand GNAME7132(G7132,G1477,G21537);
  nand GNAME7133(G7133,G29,G2263);
  nand GNAME7134(G7134,G7132,G7133);
  nand GNAME7135(G7135,G1477,G21538);
  nand GNAME7136(G7136,G30,G2263);
  nand GNAME7137(G7137,G7135,G7136);
  nand GNAME7138(G7138,G1477,G21539);
  nand GNAME7139(G7139,G31,G2263);
  nand GNAME7140(G7140,G7138,G7139);
  nand GNAME7141(G7141,G1477,G21540);
  nand GNAME7142(G7142,G32,G2263);
  nand GNAME7143(G7143,G7141,G7142);
  nand GNAME7144(G7144,G1485,G21541);
  nand GNAME7145(G7145,G25,G2262);
  nand GNAME7146(G7146,G7144,G7145);
  nand GNAME7147(G7147,G1485,G21542);
  nand GNAME7148(G7148,G26,G2262);
  nand GNAME7149(G7149,G7147,G7148);
  nand GNAME7150(G7150,G1485,G21543);
  nand GNAME7151(G7151,G27,G2262);
  nand GNAME7152(G7152,G7150,G7151);
  nand GNAME7153(G7153,G1485,G21544);
  nand GNAME7154(G7154,G28,G2262);
  nand GNAME7155(G7155,G7153,G7154);
  nand GNAME7156(G7156,G1485,G21545);
  nand GNAME7157(G7157,G29,G2262);
  nand GNAME7158(G7158,G7156,G7157);
  nand GNAME7159(G7159,G1485,G21546);
  nand GNAME7160(G7160,G30,G2262);
  nand GNAME7161(G7161,G7159,G7160);
  nand GNAME7162(G7162,G1485,G21547);
  nand GNAME7163(G7163,G31,G2262);
  nand GNAME7164(G7164,G7162,G7163);
  nand GNAME7165(G7165,G1485,G21548);
  nand GNAME7166(G7166,G32,G2262);
  nand GNAME7167(G7167,G7165,G7166);
  nand GNAME7168(G7168,G1493,G21549);
  nand GNAME7169(G7169,G25,G2261);
  nand GNAME7170(G7170,G7168,G7169);
  nand GNAME7171(G7171,G1493,G21550);
  nand GNAME7172(G7172,G26,G2261);
  nand GNAME7173(G7173,G7171,G7172);
  nand GNAME7174(G7174,G1493,G21551);
  nand GNAME7175(G7175,G27,G2261);
  nand GNAME7176(G7176,G7174,G7175);
  nand GNAME7177(G7177,G1493,G21552);
  nand GNAME7178(G7178,G28,G2261);
  nand GNAME7179(G7179,G7177,G7178);
  nand GNAME7180(G7180,G1493,G21553);
  nand GNAME7181(G7181,G29,G2261);
  nand GNAME7182(G7182,G7180,G7181);
  nand GNAME7183(G7183,G1493,G21554);
  nand GNAME7184(G7184,G30,G2261);
  nand GNAME7185(G7185,G7183,G7184);
  nand GNAME7186(G7186,G1493,G21555);
  nand GNAME7187(G7187,G31,G2261);
  nand GNAME7188(G7188,G7186,G7187);
  nand GNAME7189(G7189,G1493,G21556);
  nand GNAME7190(G7190,G32,G2261);
  nand GNAME7191(G7191,G7189,G7190);
  nand GNAME7192(G7192,G2252,G7813,G1283,G2325);
  or GNAME7193(G7193,G7289,G2252);
  nand GNAME7194(G7194,G4127,G2579);
  nand GNAME7195(G7195,G1252,G1240,G2528);
  or GNAME7196(G7196,G2494,G2253);
  nand GNAME7197(G7197,G4131,G2494);
  nand GNAME7198(G7198,G2545,G2596,G2579);
  nand GNAME7199(G7199,G1238,G1240);
  nand GNAME7200(G7200,G683,G2511);
  nand GNAME7201(G7201,G1248,G4129);
  nand GNAME7202(G7202,G4117,G21558);
  nand GNAME7203(G7203,G1213,G4116,G7207);
  not GNAME7204(G7204,G1741);
  or GNAME7205(G7205,G1213,G2252);
  nand GNAME7206(G7206,G2252,G4145);
  nand GNAME7207(G7207,G1248,G21559);
  nand GNAME7208(G7208,G1212,G2511);
  nand GNAME7209(G7209,G7207,G7208);
  nand GNAME7210(G7210,G2340,G21559);
  nand GNAME7211(G7211,G1212,G2254);
  or GNAME7212(G7212,G1212,G2252);
  nand GNAME7213(G7213,G2252,G4157);
  or GNAME7214(G7214,G1211,G2252);
  nand GNAME7215(G7215,G2252,G4172);
  or GNAME7216(G7216,G1210,G2252);
  nand GNAME7217(G7217,G2252,G4183);
  or GNAME7218(G7218,G1285,G1532);
  nand GNAME7219(G7219,G1532,G4199);
  nand GNAME7220(G7220,G1586,G21790);
  nand GNAME7221(G7221,G2330,G1199,G1207);
  nand GNAME7222(G7222,G1586,G21791);
  nand GNAME7223(G7223,G2330,G6751,G1199,G1207);
  nand GNAME7224(G7224,G1586,G21793);
  nand GNAME7225(G7225,G21758,G2330);
  nand GNAME7226(G7226,G2313,G21794);
  or GNAME7227(G7227,G21803,G2313);
  nand GNAME7228(G7228,G21797,G6772);
  nand GNAME7229(G7229,G1736,G34);
  nand GNAME7230(G7230,G21798,G2255);
  or GNAME7231(G7231,G2255,G5214);
  nand GNAME7232(G7232,G2313,G21799);
  or GNAME7233(G7233,G21801,G2313);
  nand GNAME7234(G7234,G2313,G21800);
  nand GNAME7235(G7235,G1195,G21804);
  nand GNAME7236(G7236,G21803,G2256);
  or GNAME7237(G7237,G2256,G5219);
  nand GNAME7238(G7238,G21804,G2256);
  or GNAME7239(G7239,G1296,G2256);
  nand GNAME7240(G7240,G1211,G21558);
  nand GNAME7241(G7241,G21560,G1228);
  nand GNAME7242(G7242,G1211,G21559);
  nand GNAME7243(G7243,G1212,G21560);
  not GNAME7244(G7244,G1731);
  or GNAME7245(G7245,G21795,G1212);
  nand GNAME7246(G7246,G21795,G6787,G2259);
  or GNAME7247(G7247,G21795,G1211);
  nand GNAME7248(G7248,G21795,G6787,G1727);
  or GNAME7249(G7249,G21795,G1210);
  nand GNAME7250(G7250,G4179,G21795);
  nand GNAME7251(G7251,G2257,G2325,G7813);
  or GNAME7252(G7252,G7289,G2257);
  or GNAME7253(G7253,G1213,G2257);
  nand GNAME7254(G7254,G2257,G4142);
  or GNAME7255(G7255,G1212,G2257);
  nand GNAME7256(G7256,G2257,G4153);
  or GNAME7257(G7257,G1211,G2257);
  nand GNAME7258(G7258,G2257,G4168);
  or GNAME7259(G7259,G1210,G2257);
  nand GNAME7260(G7260,G2257,G4178);
  nand GNAME7261(G7261,G1272,G21757);
  nand GNAME7262(G7262,G21427,G21598);
  nand GNAME7263(G7263,G2511,G21597);
  nand GNAME7264(G7264,G1248,G5628);
  nand GNAME7265(G7265,G2511,G21596);
  nand GNAME7266(G7266,G1248,G5645);
  nand GNAME7267(G7267,G2511,G21595);
  nand GNAME7268(G7268,G1248,G5662);
  nand GNAME7269(G7269,G2511,G21594);
  nand GNAME7270(G7270,G1248,G5679);
  nand GNAME7271(G7271,G2511,G21593);
  nand GNAME7272(G7272,G1248,G5696);
  nand GNAME7273(G7273,G2511,G21592);
  nand GNAME7274(G7274,G1248,G5713);
  nand GNAME7275(G7275,G2511,G21591);
  nand GNAME7276(G7276,G1248,G5730);
  nand GNAME7277(G7277,G2511,G21590);
  nand GNAME7278(G7278,G1248,G5747);
  nand GNAME7279(G7279,G1249,G1518);
  nand GNAME7280(G7280,G2528,G2562);
  nand GNAME7281(G7281,G1239,G1249);
  nand GNAME7282(G7282,G2562,G1242,G1192);
  nand GNAME7283(G7283,G1239,G2545);
  nand GNAME7284(G7284,G1238,G2562);
  nand GNAME7285(G7285,G21425,G21560);
  nand GNAME7286(G7286,G1208,G6716);
  nand GNAME7287(G7287,G21425,G21561);
  nand GNAME7288(G7288,G1208,G6719);
  not GNAME7289(G7289,G21557);
  not GNAME7290(G7290,G1267);
  not GNAME7291(G7291,G1318);
  not GNAME7292(G7292,G21798);
  not GNAME7293(G7293,G21562);
  not GNAME7294(G7294,G1659);
  nand GNAME7295(G7295,G7296,G21567);
  not GNAME7296(G7296,G21568);
  nand GNAME7297(G7297,G7295,G684);
  not GNAME7298(G7298,G8723);
  nand GNAME7299(G7299,G8726,G8724);
  or GNAME7300(G7300,G8724,G8726);
  nand GNAME7301(G7301,G8725,G8795);
  or GNAME7302(G7302,G8795,G8725);
  nand GNAME7303(G7303,G8729,G8728);
  or GNAME7304(G7304,G8728,G8729);
  nand GNAME7305(G7305,G8727,G8794);
  or GNAME7306(G7306,G8794,G8727);
  nand GNAME7307(G7307,G8732,G8731);
  or GNAME7308(G7308,G8731,G8732);
  nand GNAME7309(G7309,G8730,G8793);
  or GNAME7310(G7310,G8793,G8730);
  or GNAME7311(G7311,G8733,G8778);
  nand GNAME7312(G7312,G8733,G8778);
  or GNAME7313(G7313,G756,G8734);
  nand GNAME7314(G7314,G8734,G756);
  or GNAME7315(G7315,G7317,G8792);
  nand GNAME7316(G7316,G8792,G7319,G7318);
  and GNAME7317(G7317,G7319,G7318);
  nand GNAME7318(G7318,G8736,G731);
  nand GNAME7319(G7319,G8735,G755);
  not GNAME7320(G7320,G590);
  not GNAME7321(G7321,G581);
  not GNAME7322(G7322,G588);
  not GNAME7323(G7323,G579);
  not GNAME7324(G7324,G586);
  not GNAME7325(G7325,G585);
  nand GNAME7326(G7326,G7353,G7354);
  not GNAME7327(G7327,G583);
  nand GNAME7328(G7328,G7320,G582);
  nand GNAME7329(G7329,G591,G7327,G7328);
  or GNAME7330(G7330,G582,G7320);
  nand GNAME7331(G7331,G7321,G589);
  nand GNAME7332(G7332,G7331,G7329,G7330);
  or GNAME7333(G7333,G589,G7321);
  nand GNAME7334(G7334,G7322,G580);
  nand GNAME7335(G7335,G7334,G7332,G7333);
  or GNAME7336(G7336,G580,G7322);
  nand GNAME7337(G7337,G7323,G587);
  nand GNAME7338(G7338,G7337,G7335,G7336);
  or GNAME7339(G7339,G587,G7323);
  nand GNAME7340(G7340,G7324,G578);
  nand GNAME7341(G7341,G7340,G7338,G7339);
  or GNAME7342(G7342,G578,G7324);
  or GNAME7343(G7343,G578,G7325);
  nand GNAME7344(G7344,G7343,G7341,G7342);
  nand GNAME7345(G7345,G7325,G578);
  and GNAME7346(G7346,G7345,G7344);
  nand GNAME7347(G7347,G576,G584);
  or GNAME7348(G7348,G584,G7346);
  and GNAME7349(G7349,G7347,G7348);
  or GNAME7350(G7350,G576,G584);
  or GNAME7351(G7351,G7346,G7355);
  nand GNAME7352(G7352,G7350,G7351);
  or GNAME7353(G7353,G577,G7349);
  nand GNAME7354(G7354,G7352,G577);
  not GNAME7355(G7355,G584);
  not GNAME7356(G7356,G7436);
  nand GNAME7357(G7357,G7581,G7436);
  not GNAME7358(G7358,G7435);
  nand GNAME7359(G7359,G7580,G7435);
  not GNAME7360(G7360,G7434);
  nand GNAME7361(G7361,G7579,G7434);
  not GNAME7362(G7362,G7433);
  nand GNAME7363(G7363,G7578,G7433);
  not GNAME7364(G7364,G7432);
  nand GNAME7365(G7365,G7577,G7432);
  not GNAME7366(G7366,G7431);
  nand GNAME7367(G7367,G7576,G7431);
  not GNAME7368(G7368,G7430);
  nand GNAME7369(G7369,G7575,G7430);
  not GNAME7370(G7370,G7429);
  nand GNAME7371(G7371,G7574,G7429);
  not GNAME7372(G7372,G7428);
  nand GNAME7373(G7373,G7573,G7428);
  not GNAME7374(G7374,G7427);
  nand GNAME7375(G7375,G7572,G7427);
  not GNAME7376(G7376,G7426);
  nand GNAME7377(G7377,G7571,G7426);
  not GNAME7378(G7378,G7425);
  nand GNAME7379(G7379,G7570,G7425);
  not GNAME7380(G7380,G7424);
  nand GNAME7381(G7381,G7569,G7424);
  not GNAME7382(G7382,G7423);
  nand GNAME7383(G7383,G7568,G7423);
  nand GNAME7384(G7384,G7416,G7418);
  not GNAME7385(G7385,G7418);
  not GNAME7386(G7386,G7422);
  nand GNAME7387(G7387,G7538,G7422);
  not GNAME7388(G7388,G7391);
  nand GNAME7389(G7389,G7532,G7391);
  not GNAME7390(G7390,G7531);
  nand GNAME7391(G7391,G7622,G7623);
  and GNAME7392(G7392,G7420,G7390);
  and GNAME7393(G7393,G7392,G7391);
  and GNAME7394(G7394,G7707,G7415);
  and GNAME7395(G7395,G7418,G7394);
  and GNAME7396(G7396,G7520,G7423);
  and GNAME7397(G7397,G7396,G7424);
  and GNAME7398(G7398,G7397,G7425);
  and GNAME7399(G7399,G7398,G7426);
  and GNAME7400(G7400,G7399,G7427);
  and GNAME7401(G7401,G7400,G7428);
  and GNAME7402(G7402,G7401,G7429);
  and GNAME7403(G7403,G7402,G7430);
  and GNAME7404(G7404,G7403,G7431);
  and GNAME7405(G7405,G7404,G7432);
  and GNAME7406(G7406,G7405,G7433);
  and GNAME7407(G7407,G7406,G7434);
  and GNAME7408(G7408,G7407,G7435);
  nand GNAME7409(G7409,G7410,G7420);
  not GNAME7410(G7410,G7460);
  nand GNAME7411(G7411,G7412,G7460);
  not GNAME7412(G7412,G7420);
  nand GNAME7413(G7413,G7634,G7458);
  and GNAME7414(G7414,G7635,G7636);
  not GNAME7415(G7415,G7539);
  not GNAME7416(G7416,G7451);
  nand GNAME7417(G7417,G7385,G7451);
  nand GNAME7418(G7418,G7607,G7608);
  and GNAME7419(G7419,G7609,G7610);
  nand GNAME7420(G7420,G7613,G7614);
  and GNAME7421(G7421,G7615,G7616);
  nand GNAME7422(G7422,G7611,G7612);
  nand GNAME7423(G7423,G7655,G7656);
  nand GNAME7424(G7424,G7657,G7658);
  nand GNAME7425(G7425,G7659,G7660);
  nand GNAME7426(G7426,G7661,G7662);
  nand GNAME7427(G7427,G7663,G7664);
  nand GNAME7428(G7428,G7665,G7666);
  nand GNAME7429(G7429,G7667,G7668);
  nand GNAME7430(G7430,G7669,G7670);
  nand GNAME7431(G7431,G7671,G7672);
  nand GNAME7432(G7432,G7673,G7674);
  nand GNAME7433(G7433,G7675,G7676);
  nand GNAME7434(G7434,G7677,G7678);
  nand GNAME7435(G7435,G7679,G7680);
  nand GNAME7436(G7436,G7681,G7682);
  and GNAME7437(G7437,G7595,G7596);
  and GNAME7438(G7438,G7591,G7593);
  and GNAME7439(G7439,G7587,G7588);
  and GNAME7440(G7440,G7585,G7460);
  and GNAME7441(G7441,G7710,G7584);
  and GNAME7442(G7442,G7413,G7583);
  and GNAME7443(G7443,G7409,G7411);
  and GNAME7444(G7444,G7540,G7451);
  and GNAME7445(G7445,G7384,G7417);
  not GNAME7446(G7446,G2297);
  not GNAME7447(G7447,G633);
  not GNAME7448(G7448,G632);
  not GNAME7449(G7449,G631);
  not GNAME7450(G7450,G630);
  or GNAME7451(G7451,G7419,G7539);
  not GNAME7452(G7452,G629);
  not GNAME7453(G7453,G628);
  not GNAME7454(G7454,G627);
  not GNAME7455(G7455,G626);
  not GNAME7456(G7456,G625);
  not GNAME7457(G7457,G624);
  nor GNAME7458(G7458,G7414,G7582);
  and GNAME7459(G7459,G7543,G7528);
  or GNAME7460(G7460,G7421,G7459);
  and GNAME7461(G7461,G7564,G7563);
  nor GNAME7462(G7462,G7565,G7461);
  and GNAME7463(G7463,G7589,G7537);
  or GNAME7464(G7464,G7549,G7463);
  and GNAME7465(G7465,G7619,G7620);
  and GNAME7466(G7466,G7624,G7625);
  nand GNAME7467(G7467,G7705,G7706);
  nand GNAME7468(G7468,G7626,G7627);
  nand GNAME7469(G7469,G7628,G7629);
  nand GNAME7470(G7470,G7630,G7387);
  nand GNAME7471(G7471,G7631,G7389);
  nand GNAME7472(G7472,G7683,G7357);
  nand GNAME7473(G7473,G7684,G7359);
  nand GNAME7474(G7474,G7685,G7361);
  nand GNAME7475(G7475,G7686,G7363);
  nand GNAME7476(G7476,G7687,G7365);
  nand GNAME7477(G7477,G7688,G7367);
  nand GNAME7478(G7478,G7689,G7369);
  nand GNAME7479(G7479,G7690,G7371);
  nand GNAME7480(G7480,G7691,G7373);
  nand GNAME7481(G7481,G7692,G7375);
  nand GNAME7482(G7482,G7693,G7694);
  nand GNAME7483(G7483,G7695,G7377);
  nand GNAME7484(G7484,G7696,G7379);
  nand GNAME7485(G7485,G7697,G7381);
  nand GNAME7486(G7486,G7698,G7383);
  nand GNAME7487(G7487,G7699,G7700);
  nand GNAME7488(G7488,G7701,G7702);
  nand GNAME7489(G7489,G7703,G7704);
  not GNAME7490(G7490,G614);
  not GNAME7491(G7491,G616);
  not GNAME7492(G7492,G617);
  not GNAME7493(G7493,G618);
  not GNAME7494(G7494,G620);
  not GNAME7495(G7495,G621);
  not GNAME7496(G7496,G622);
  not GNAME7497(G7497,G592);
  not GNAME7498(G7498,G593);
  not GNAME7499(G7499,G608);
  not GNAME7500(G7500,G609);
  not GNAME7501(G7501,G612);
  not GNAME7502(G7502,G613);
  not GNAME7503(G7503,G611);
  not GNAME7504(G7504,G610);
  not GNAME7505(G7505,G607);
  not GNAME7506(G7506,G606);
  not GNAME7507(G7507,G605);
  not GNAME7508(G7508,G604);
  not GNAME7509(G7509,G603);
  not GNAME7510(G7510,G602);
  not GNAME7511(G7511,G601);
  not GNAME7512(G7512,G600);
  not GNAME7513(G7513,G599);
  not GNAME7514(G7514,G598);
  not GNAME7515(G7515,G597);
  not GNAME7516(G7516,G596);
  not GNAME7517(G7517,G595);
  not GNAME7518(G7518,G594);
  nand GNAME7519(G7519,G7541,G7526);
  nand GNAME7520(G7520,G7567,G7545);
  or GNAME7521(G7521,G7462,G7546);
  nand GNAME7522(G7522,G7560,G7559);
  nand GNAME7523(G7523,G7556,G7548);
  nand GNAME7524(G7524,G7529,G7526);
  or GNAME7525(G7525,G7466,G7449);
  or GNAME7526(G7526,G7465,G7447);
  nand GNAME7527(G7527,G7448,G7617,G7618);
  nand GNAME7528(G7528,G7621,G632);
  nand GNAME7529(G7529,G7447,G7465);
  nand GNAME7530(G7530,G7543,G7528);
  nand GNAME7531(G7531,G7708,G7530);
  not GNAME7532(G7532,G7392);
  not GNAME7533(G7533,G7395);
  nand GNAME7534(G7534,G7449,G7466);
  not GNAME7535(G7535,G7552);
  nand GNAME7536(G7536,G7450,G7604,G7605);
  nand GNAME7537(G7537,G7606,G630);
  not GNAME7538(G7538,G7393);
  nand GNAME7539(G7539,G7422,G7393);
  nand GNAME7540(G7540,G7419,G7539);
  nand GNAME7541(G7541,G7529,G2297);
  not GNAME7542(G7542,G7519);
  nand GNAME7543(G7543,G7527,G7519);
  nand GNAME7544(G7544,G7457,G7637,G7638);
  nand GNAME7545(G7545,G7654,G624);
  and GNAME7546(G7546,G7653,G625);
  nand GNAME7547(G7547,G7453,G7641,G7642);
  nand GNAME7548(G7548,G7646,G628);
  and GNAME7549(G7549,G7452,G7643,G7644);
  nand GNAME7550(G7550,G7645,G629);
  nand GNAME7551(G7551,G7395,G7534);
  nand GNAME7552(G7552,G7551,G7525);
  nand GNAME7553(G7553,G7589,G7537);
  nand GNAME7554(G7554,G7709,G7553);
  nand GNAME7555(G7555,G7554,G7550);
  nand GNAME7556(G7556,G7547,G7555);
  not GNAME7557(G7557,G7523);
  nand GNAME7558(G7558,G7454,G7647,G7648);
  nand GNAME7559(G7559,G7649,G627);
  nand GNAME7560(G7560,G7523,G7558);
  not GNAME7561(G7561,G7522);
  nand GNAME7562(G7562,G7455,G7650,G7651);
  nand GNAME7563(G7563,G7652,G626);
  nand GNAME7564(G7564,G7522,G7562);
  and GNAME7565(G7565,G7456,G7639,G7640);
  not GNAME7566(G7566,G7521);
  nand GNAME7567(G7567,G7544,G7521);
  not GNAME7568(G7568,G7520);
  not GNAME7569(G7569,G7396);
  not GNAME7570(G7570,G7397);
  not GNAME7571(G7571,G7398);
  not GNAME7572(G7572,G7399);
  not GNAME7573(G7573,G7400);
  not GNAME7574(G7574,G7401);
  not GNAME7575(G7575,G7402);
  not GNAME7576(G7576,G7403);
  not GNAME7577(G7577,G7404);
  not GNAME7578(G7578,G7405);
  not GNAME7579(G7579,G7406);
  not GNAME7580(G7580,G7407);
  not GNAME7581(G7581,G7408);
  nand GNAME7582(G7582,G7408,G7436);
  nand GNAME7583(G7583,G7710,G7632,G7633);
  nand GNAME7584(G7584,G7414,G7582);
  nand GNAME7585(G7585,G7421,G7459);
  or GNAME7586(G7586,G7546,G7565);
  nand GNAME7587(G7587,G7586,G7461);
  or GNAME7588(G7588,G7546,G7711);
  nand GNAME7589(G7589,G7552,G7536);
  nand GNAME7590(G7590,G7550,G7464);
  nand GNAME7591(G7591,G7590,G7547,G7548);
  nand GNAME7592(G7592,G7547,G7548);
  nand GNAME7593(G7593,G7592,G7550,G7464);
  or GNAME7594(G7594,G7549,G7712);
  nand GNAME7595(G7595,G7594,G7463);
  or GNAME7596(G7596,G7712,G7464);
  not GNAME7597(G7597,G7524);
  nand GNAME7598(G7598,G7536,G7537);
  nand GNAME7599(G7599,G7525,G7534);
  nand GNAME7600(G7600,G7527,G7528);
  nand GNAME7601(G7601,G7544,G7545);
  nand GNAME7602(G7602,G7562,G7563);
  nand GNAME7603(G7603,G7558,G7559);
  nand GNAME7604(G7604,G7490,G2297);
  nand GNAME7605(G7605,G7446,G614);
  nand GNAME7606(G7606,G7604,G7605);
  nand GNAME7607(G7607,G7491,G2297);
  nand GNAME7608(G7608,G7446,G616);
  nand GNAME7609(G7609,G7492,G2297);
  nand GNAME7610(G7610,G7446,G617);
  nand GNAME7611(G7611,G7493,G2297);
  nand GNAME7612(G7612,G7446,G618);
  nand GNAME7613(G7613,G7494,G2297);
  nand GNAME7614(G7614,G7446,G620);
  nand GNAME7615(G7615,G7495,G2297);
  nand GNAME7616(G7616,G7446,G621);
  nand GNAME7617(G7617,G7496,G2297);
  nand GNAME7618(G7618,G7446,G622);
  or GNAME7619(G7619,G623,G7446);
  nand GNAME7620(G7620,G7446,G623);
  nand GNAME7621(G7621,G7617,G7618);
  or GNAME7622(G7622,G619,G7446);
  nand GNAME7623(G7623,G7446,G619);
  or GNAME7624(G7624,G615,G7446);
  nand GNAME7625(G7625,G7446,G615);
  nand GNAME7626(G7626,G7552,G7598);
  nand GNAME7627(G7627,G7535,G7536,G7537);
  nand GNAME7628(G7628,G7395,G7599);
  nand GNAME7629(G7629,G7533,G7525,G7534);
  nand GNAME7630(G7630,G7393,G7386);
  nand GNAME7631(G7631,G7392,G7388);
  nand GNAME7632(G7632,G7497,G2297);
  nand GNAME7633(G7633,G7446,G592);
  nand GNAME7634(G7634,G7632,G7633);
  nand GNAME7635(G7635,G7498,G2297);
  nand GNAME7636(G7636,G7446,G593);
  nand GNAME7637(G7637,G7499,G2297);
  nand GNAME7638(G7638,G7446,G608);
  nand GNAME7639(G7639,G7500,G2297);
  nand GNAME7640(G7640,G7446,G609);
  nand GNAME7641(G7641,G7501,G2297);
  nand GNAME7642(G7642,G7446,G612);
  nand GNAME7643(G7643,G7502,G2297);
  nand GNAME7644(G7644,G7446,G613);
  nand GNAME7645(G7645,G7643,G7644);
  nand GNAME7646(G7646,G7641,G7642);
  nand GNAME7647(G7647,G7503,G2297);
  nand GNAME7648(G7648,G7446,G611);
  nand GNAME7649(G7649,G7647,G7648);
  nand GNAME7650(G7650,G7504,G2297);
  nand GNAME7651(G7651,G7446,G610);
  nand GNAME7652(G7652,G7650,G7651);
  nand GNAME7653(G7653,G7639,G7640);
  nand GNAME7654(G7654,G7637,G7638);
  nand GNAME7655(G7655,G7505,G2297);
  nand GNAME7656(G7656,G7446,G607);
  nand GNAME7657(G7657,G7506,G2297);
  nand GNAME7658(G7658,G7446,G606);
  nand GNAME7659(G7659,G7507,G2297);
  nand GNAME7660(G7660,G7446,G605);
  nand GNAME7661(G7661,G7508,G2297);
  nand GNAME7662(G7662,G7446,G604);
  nand GNAME7663(G7663,G7509,G2297);
  nand GNAME7664(G7664,G7446,G603);
  nand GNAME7665(G7665,G7510,G2297);
  nand GNAME7666(G7666,G7446,G602);
  nand GNAME7667(G7667,G7511,G2297);
  nand GNAME7668(G7668,G7446,G601);
  nand GNAME7669(G7669,G7512,G2297);
  nand GNAME7670(G7670,G7446,G600);
  nand GNAME7671(G7671,G7513,G2297);
  nand GNAME7672(G7672,G7446,G599);
  nand GNAME7673(G7673,G7514,G2297);
  nand GNAME7674(G7674,G7446,G598);
  nand GNAME7675(G7675,G7515,G2297);
  nand GNAME7676(G7676,G7446,G597);
  nand GNAME7677(G7677,G7516,G2297);
  nand GNAME7678(G7678,G7446,G596);
  nand GNAME7679(G7679,G7517,G2297);
  nand GNAME7680(G7680,G7446,G595);
  nand GNAME7681(G7681,G7518,G2297);
  nand GNAME7682(G7682,G7446,G594);
  nand GNAME7683(G7683,G7408,G7356);
  nand GNAME7684(G7684,G7407,G7358);
  nand GNAME7685(G7685,G7406,G7360);
  nand GNAME7686(G7686,G7405,G7362);
  nand GNAME7687(G7687,G7404,G7364);
  nand GNAME7688(G7688,G7403,G7366);
  nand GNAME7689(G7689,G7402,G7368);
  nand GNAME7690(G7690,G7401,G7370);
  nand GNAME7691(G7691,G7400,G7372);
  nand GNAME7692(G7692,G7399,G7374);
  nand GNAME7693(G7693,G7519,G7600);
  nand GNAME7694(G7694,G7542,G7527,G7528);
  nand GNAME7695(G7695,G7398,G7376);
  nand GNAME7696(G7696,G7397,G7378);
  nand GNAME7697(G7697,G7396,G7380);
  nand GNAME7698(G7698,G7520,G7382);
  nand GNAME7699(G7699,G7521,G7601);
  nand GNAME7700(G7700,G7566,G7544,G7545);
  nand GNAME7701(G7701,G7522,G7602);
  nand GNAME7702(G7702,G7561,G7562,G7563);
  nand GNAME7703(G7703,G7523,G7603);
  nand GNAME7704(G7704,G7557,G7558,G7559);
  nand GNAME7705(G7705,G7524,G2297);
  nand GNAME7706(G7706,G7446,G7597);
  not GNAME7707(G7707,G7419);
  not GNAME7708(G7708,G7421);
  not GNAME7709(G7709,G7549);
  not GNAME7710(G7710,G7458);
  not GNAME7711(G7711,G7462);
  not GNAME7712(G7712,G7550);
  not GNAME7713(G7713,G561);
  not GNAME7714(G7714,G566);
  not GNAME7715(G7715,G560);
  not GNAME7716(G7716,G562);
  not GNAME7717(G7717,G567);
  not GNAME7718(G7718,G564);
  not GNAME7719(G7719,G565);
  not GNAME7720(G7720,G563);
  and GNAME7721(G7721,G7839,G7772);
  and GNAME7722(G7722,G8097,G7760);
  and GNAME7723(G7723,G7766,G7722);
  and GNAME7724(G7724,G7723,G7761);
  and GNAME7725(G7725,G7753,G7804);
  and GNAME7726(G7726,G7864,G7750);
  and GNAME7727(G7727,G7726,G7747);
  and GNAME7728(G7728,G7727,G7744);
  and GNAME7729(G7729,G7728,G7741);
  and GNAME7730(G7730,G7729,G7738);
  nand GNAME7731(G7731,G8015,G7801);
  and GNAME7732(G7732,G8016,G8017);
  not GNAME7733(G7733,G7735);
  nand GNAME7734(G7734,G7959,G7735);
  nand GNAME7735(G7735,G8064,G8065);
  not GNAME7736(G7736,G7738);
  nand GNAME7737(G7737,G7958,G7738);
  nand GNAME7738(G7738,G8062,G8063);
  not GNAME7739(G7739,G7741);
  nand GNAME7740(G7740,G7957,G7741);
  nand GNAME7741(G7741,G8060,G8061);
  not GNAME7742(G7742,G7744);
  nand GNAME7743(G7743,G7956,G7744);
  nand GNAME7744(G7744,G8058,G8059);
  not GNAME7745(G7745,G7747);
  nand GNAME7746(G7746,G7955,G7747);
  nand GNAME7747(G7747,G8056,G8057);
  not GNAME7748(G7748,G7750);
  nand GNAME7749(G7749,G7954,G7750);
  nand GNAME7750(G7750,G8054,G8055);
  not GNAME7751(G7751,G7753);
  nand GNAME7752(G7752,G7921,G7753);
  nand GNAME7753(G7753,G8018,G8019);
  and GNAME7754(G7754,G8020,G8021);
  not GNAME7755(G7755,G7757);
  nand GNAME7756(G7756,G7919,G7757);
  nand GNAME7757(G7757,G8028,G8029);
  not GNAME7758(G7758,G7761);
  nand GNAME7759(G7759,G7918,G7761);
  not GNAME7760(G7760,G7967);
  nand GNAME7761(G7761,G8026,G8027);
  nand GNAME7762(G7762,G7763,G7766);
  not GNAME7763(G7763,G7805);
  nand GNAME7764(G7764,G7765,G7805);
  not GNAME7765(G7765,G7766);
  nand GNAME7766(G7766,G8022,G8023);
  and GNAME7767(G7767,G8024,G8025);
  not GNAME7768(G7768,G7770);
  nand GNAME7769(G7769,G7900,G7770);
  nand GNAME7770(G7770,G7981,G7982);
  nand GNAME7771(G7771,G7899,G7772);
  not GNAME7772(G7772,G7808);
  and GNAME7773(G7773,G7968,G7805);
  and GNAME7774(G7774,G7762,G7764);
  and GNAME7775(G7775,G7966,G7921);
  and GNAME7776(G7776,G7964,G7965);
  and GNAME7777(G7777,G8099,G7962);
  and GNAME7778(G7778,G7731,G7961);
  and GNAME7779(G7779,G7915,G7917);
  and GNAME7780(G7780,G7909,G7910);
  and GNAME7781(G7781,G7905,G7907);
  not GNAME7782(G7782,G1278);
  not GNAME7783(G7783,G681);
  not GNAME7784(G7784,G680);
  not GNAME7785(G7785,G679);
  not GNAME7786(G7786,G678);
  not GNAME7787(G7787,G677);
  not GNAME7788(G7788,G676);
  not GNAME7789(G7789,G675);
  not GNAME7790(G7790,G674);
  and GNAME7791(G7791,G7903,G7881);
  or GNAME7792(G7792,G7878,G7791);
  not GNAME7793(G7793,G673);
  not GNAME7794(G7794,G672);
  not GNAME7795(G7795,G671);
  not GNAME7796(G7796,G670);
  not GNAME7797(G7797,G669);
  not GNAME7798(G7798,G668);
  not GNAME7799(G7799,G667);
  not GNAME7800(G7800,G666);
  nor GNAME7801(G7801,G7732,G7960);
  and GNAME7802(G7802,G7913,G7887);
  or GNAME7803(G7803,G7884,G7802);
  nor GNAME7804(G7804,G7754,G7920);
  or GNAME7805(G7805,G7767,G7967);
  and GNAME7806(G7806,G7995,G7996);
  and GNAME7807(G7807,G8000,G8001);
  and GNAME7808(G7808,G8005,G8006);
  nand GNAME7809(G7809,G8093,G8094);
  nand GNAME7810(G7810,G8007,G7769);
  nand GNAME7811(G7811,G8008,G7771);
  nand GNAME7812(G7812,G8009,G8010);
  nand GNAME7813(G7813,G8011,G8012);
  nand GNAME7814(G7814,G8066,G7734);
  nand GNAME7815(G7815,G8067,G7737);
  nand GNAME7816(G7816,G8068,G7740);
  nand GNAME7817(G7817,G8069,G7743);
  nand GNAME7818(G7818,G8070,G7746);
  nand GNAME7819(G7819,G8071,G7749);
  nand GNAME7820(G7820,G8072,G8073);
  nand GNAME7821(G7821,G8074,G8075);
  nand GNAME7822(G7822,G8076,G8077);
  nand GNAME7823(G7823,G8078,G8079);
  nand GNAME7824(G7824,G8080,G8081);
  nand GNAME7825(G7825,G8082,G8083);
  nand GNAME7826(G7826,G8084,G8085);
  nand GNAME7827(G7827,G8086,G8087);
  nand GNAME7828(G7828,G8088,G8089);
  nand GNAME7829(G7829,G8090,G7752);
  nand GNAME7830(G7830,G8091,G7756);
  nand GNAME7831(G7831,G8092,G7759);
  not GNAME7832(G7832,G656);
  not GNAME7833(G7833,G658);
  not GNAME7834(G7834,G659);
  not GNAME7835(G7835,G660);
  not GNAME7836(G7836,G662);
  not GNAME7837(G7837,G663);
  not GNAME7838(G7838,G664);
  nand GNAME7839(G7839,G7898,G7877);
  nand GNAME7840(G7840,G7901,G7875);
  nand GNAME7841(G7841,G7892,G7883);
  not GNAME7842(G7842,G634);
  not GNAME7843(G7843,G635);
  not GNAME7844(G7844,G650);
  not GNAME7845(G7845,G651);
  not GNAME7846(G7846,G654);
  not GNAME7847(G7847,G655);
  not GNAME7848(G7848,G653);
  not GNAME7849(G7849,G652);
  not GNAME7850(G7850,G649);
  not GNAME7851(G7851,G648);
  not GNAME7852(G7852,G647);
  not GNAME7853(G7853,G646);
  not GNAME7854(G7854,G645);
  not GNAME7855(G7855,G644);
  not GNAME7856(G7856,G643);
  not GNAME7857(G7857,G642);
  not GNAME7858(G7858,G641);
  not GNAME7859(G7859,G640);
  not GNAME7860(G7860,G639);
  not GNAME7861(G7861,G638);
  not GNAME7862(G7862,G637);
  not GNAME7863(G7863,G636);
  nand GNAME7864(G7864,G7953,G7952);
  nand GNAME7865(G7865,G7949,G7948);
  nand GNAME7866(G7866,G7945,G7944);
  nand GNAME7867(G7867,G7941,G7940);
  nand GNAME7868(G7868,G7937,G7936);
  nand GNAME7869(G7869,G7911,G7874);
  nand GNAME7870(G7870,G7933,G7932);
  nand GNAME7871(G7871,G7929,G7928);
  nand GNAME7872(G7872,G7925,G7924);
  nand GNAME7873(G7873,G7888,G7874);
  or GNAME7874(G7874,G7806,G7783);
  or GNAME7875(G7875,G7807,G7787);
  nand GNAME7876(G7876,G7790,G7983,G7984);
  nand GNAME7877(G7877,G8004,G674);
  and GNAME7878(G7878,G7789,G7985,G7986);
  nand GNAME7879(G7879,G8003,G675);
  nand GNAME7880(G7880,G7788,G7987,G7988);
  nand GNAME7881(G7881,G8002,G676);
  nand GNAME7882(G7882,G7786,G7989,G7990);
  nand GNAME7883(G7883,G7999,G678);
  and GNAME7884(G7884,G7785,G7991,G7992);
  nand GNAME7885(G7885,G7998,G679);
  nand GNAME7886(G7886,G7784,G7993,G7994);
  nand GNAME7887(G7887,G7997,G680);
  nand GNAME7888(G7888,G7783,G7806);
  nand GNAME7889(G7889,G7913,G7887);
  nand GNAME7890(G7890,G8096,G7889);
  nand GNAME7891(G7891,G7890,G7885);
  nand GNAME7892(G7892,G7882,G7891);
  not GNAME7893(G7893,G7841);
  nand GNAME7894(G7894,G7787,G7807);
  nand GNAME7895(G7895,G7903,G7881);
  nand GNAME7896(G7896,G8095,G7895);
  nand GNAME7897(G7897,G7896,G7879);
  nand GNAME7898(G7898,G7876,G7897);
  not GNAME7899(G7899,G7839);
  not GNAME7900(G7900,G7721);
  nand GNAME7901(G7901,G7841,G7894);
  not GNAME7902(G7902,G7840);
  nand GNAME7903(G7903,G7880,G7840);
  nand GNAME7904(G7904,G7879,G7792);
  nand GNAME7905(G7905,G7904,G7876,G7877);
  nand GNAME7906(G7906,G7876,G7877);
  nand GNAME7907(G7907,G7906,G7879,G7792);
  or GNAME7908(G7908,G7878,G8098);
  nand GNAME7909(G7909,G7908,G7791);
  or GNAME7910(G7910,G8098,G7792);
  nand GNAME7911(G7911,G7888,G1278);
  not GNAME7912(G7912,G7869);
  nand GNAME7913(G7913,G7886,G7869);
  nand GNAME7914(G7914,G7885,G7803);
  nand GNAME7915(G7915,G7914,G7882,G7883);
  nand GNAME7916(G7916,G7882,G7883);
  nand GNAME7917(G7917,G7916,G7885,G7803);
  not GNAME7918(G7918,G7723);
  not GNAME7919(G7919,G7724);
  nand GNAME7920(G7920,G7724,G7757);
  not GNAME7921(G7921,G7804);
  not GNAME7922(G7922,G7725);
  nand GNAME7923(G7923,G7793,G8030,G8031);
  nand GNAME7924(G7924,G8032,G673);
  nand GNAME7925(G7925,G7725,G7923);
  not GNAME7926(G7926,G7872);
  nand GNAME7927(G7927,G7794,G8033,G8034);
  nand GNAME7928(G7928,G8035,G672);
  nand GNAME7929(G7929,G7872,G7927);
  not GNAME7930(G7930,G7871);
  nand GNAME7931(G7931,G7795,G8036,G8037);
  nand GNAME7932(G7932,G8038,G671);
  nand GNAME7933(G7933,G7871,G7931);
  not GNAME7934(G7934,G7870);
  nand GNAME7935(G7935,G7796,G8039,G8040);
  nand GNAME7936(G7936,G8041,G670);
  nand GNAME7937(G7937,G7870,G7935);
  not GNAME7938(G7938,G7868);
  nand GNAME7939(G7939,G7797,G8042,G8043);
  nand GNAME7940(G7940,G8044,G669);
  nand GNAME7941(G7941,G7868,G7939);
  not GNAME7942(G7942,G7867);
  nand GNAME7943(G7943,G7798,G8045,G8046);
  nand GNAME7944(G7944,G8047,G668);
  nand GNAME7945(G7945,G7867,G7943);
  not GNAME7946(G7946,G7866);
  nand GNAME7947(G7947,G7799,G8048,G8049);
  nand GNAME7948(G7948,G8050,G667);
  nand GNAME7949(G7949,G7866,G7947);
  not GNAME7950(G7950,G7865);
  nand GNAME7951(G7951,G7800,G8051,G8052);
  nand GNAME7952(G7952,G8053,G666);
  nand GNAME7953(G7953,G7865,G7951);
  not GNAME7954(G7954,G7864);
  not GNAME7955(G7955,G7726);
  not GNAME7956(G7956,G7727);
  not GNAME7957(G7957,G7728);
  not GNAME7958(G7958,G7729);
  not GNAME7959(G7959,G7730);
  nand GNAME7960(G7960,G7730,G7735);
  nand GNAME7961(G7961,G8099,G8013,G8014);
  nand GNAME7962(G7962,G7732,G7960);
  or GNAME7963(G7963,G7884,G8100);
  nand GNAME7964(G7964,G7963,G7802);
  or GNAME7965(G7965,G8100,G7803);
  nand GNAME7966(G7966,G7754,G7920);
  nand GNAME7967(G7967,G7721,G7770);
  nand GNAME7968(G7968,G7767,G7967);
  not GNAME7969(G7969,G7873);
  nand GNAME7970(G7970,G7880,G7881);
  nand GNAME7971(G7971,G7875,G7894);
  nand GNAME7972(G7972,G7951,G7952);
  nand GNAME7973(G7973,G7947,G7948);
  nand GNAME7974(G7974,G7943,G7944);
  nand GNAME7975(G7975,G7939,G7940);
  nand GNAME7976(G7976,G7886,G7887);
  nand GNAME7977(G7977,G7935,G7936);
  nand GNAME7978(G7978,G7931,G7932);
  nand GNAME7979(G7979,G7927,G7928);
  nand GNAME7980(G7980,G7923,G7924);
  nand GNAME7981(G7981,G7832,G1278);
  nand GNAME7982(G7982,G7782,G656);
  nand GNAME7983(G7983,G7833,G1278);
  nand GNAME7984(G7984,G7782,G658);
  nand GNAME7985(G7985,G7834,G1278);
  nand GNAME7986(G7986,G7782,G659);
  nand GNAME7987(G7987,G7835,G1278);
  nand GNAME7988(G7988,G7782,G660);
  nand GNAME7989(G7989,G7836,G1278);
  nand GNAME7990(G7990,G7782,G662);
  nand GNAME7991(G7991,G7837,G1278);
  nand GNAME7992(G7992,G7782,G663);
  nand GNAME7993(G7993,G7838,G1278);
  nand GNAME7994(G7994,G7782,G664);
  or GNAME7995(G7995,G665,G7782);
  nand GNAME7996(G7996,G7782,G665);
  nand GNAME7997(G7997,G7993,G7994);
  nand GNAME7998(G7998,G7991,G7992);
  nand GNAME7999(G7999,G7989,G7990);
  or GNAME8000(G8000,G661,G7782);
  nand GNAME8001(G8001,G7782,G661);
  nand GNAME8002(G8002,G7987,G7988);
  nand GNAME8003(G8003,G7985,G7986);
  nand GNAME8004(G8004,G7983,G7984);
  or GNAME8005(G8005,G657,G7782);
  nand GNAME8006(G8006,G7782,G657);
  nand GNAME8007(G8007,G7721,G7768);
  nand GNAME8008(G8008,G7839,G7808);
  nand GNAME8009(G8009,G7840,G7970);
  nand GNAME8010(G8010,G7902,G7880,G7881);
  nand GNAME8011(G8011,G7841,G7971);
  nand GNAME8012(G8012,G7893,G7875,G7894);
  nand GNAME8013(G8013,G7842,G1278);
  nand GNAME8014(G8014,G7782,G634);
  nand GNAME8015(G8015,G8013,G8014);
  nand GNAME8016(G8016,G7843,G1278);
  nand GNAME8017(G8017,G7782,G635);
  nand GNAME8018(G8018,G7844,G1278);
  nand GNAME8019(G8019,G7782,G650);
  nand GNAME8020(G8020,G7845,G1278);
  nand GNAME8021(G8021,G7782,G651);
  nand GNAME8022(G8022,G7846,G1278);
  nand GNAME8023(G8023,G7782,G654);
  nand GNAME8024(G8024,G7847,G1278);
  nand GNAME8025(G8025,G7782,G655);
  nand GNAME8026(G8026,G7848,G1278);
  nand GNAME8027(G8027,G7782,G653);
  nand GNAME8028(G8028,G7849,G1278);
  nand GNAME8029(G8029,G7782,G652);
  nand GNAME8030(G8030,G7850,G1278);
  nand GNAME8031(G8031,G7782,G649);
  nand GNAME8032(G8032,G8030,G8031);
  nand GNAME8033(G8033,G7851,G1278);
  nand GNAME8034(G8034,G7782,G648);
  nand GNAME8035(G8035,G8033,G8034);
  nand GNAME8036(G8036,G7852,G1278);
  nand GNAME8037(G8037,G7782,G647);
  nand GNAME8038(G8038,G8036,G8037);
  nand GNAME8039(G8039,G7853,G1278);
  nand GNAME8040(G8040,G7782,G646);
  nand GNAME8041(G8041,G8039,G8040);
  nand GNAME8042(G8042,G7854,G1278);
  nand GNAME8043(G8043,G7782,G645);
  nand GNAME8044(G8044,G8042,G8043);
  nand GNAME8045(G8045,G7855,G1278);
  nand GNAME8046(G8046,G7782,G644);
  nand GNAME8047(G8047,G8045,G8046);
  nand GNAME8048(G8048,G7856,G1278);
  nand GNAME8049(G8049,G7782,G643);
  nand GNAME8050(G8050,G8048,G8049);
  nand GNAME8051(G8051,G7857,G1278);
  nand GNAME8052(G8052,G7782,G642);
  nand GNAME8053(G8053,G8051,G8052);
  nand GNAME8054(G8054,G7858,G1278);
  nand GNAME8055(G8055,G7782,G641);
  nand GNAME8056(G8056,G7859,G1278);
  nand GNAME8057(G8057,G7782,G640);
  nand GNAME8058(G8058,G7860,G1278);
  nand GNAME8059(G8059,G7782,G639);
  nand GNAME8060(G8060,G7861,G1278);
  nand GNAME8061(G8061,G7782,G638);
  nand GNAME8062(G8062,G7862,G1278);
  nand GNAME8063(G8063,G7782,G637);
  nand GNAME8064(G8064,G7863,G1278);
  nand GNAME8065(G8065,G7782,G636);
  nand GNAME8066(G8066,G7730,G7733);
  nand GNAME8067(G8067,G7729,G7736);
  nand GNAME8068(G8068,G7728,G7739);
  nand GNAME8069(G8069,G7727,G7742);
  nand GNAME8070(G8070,G7726,G7745);
  nand GNAME8071(G8071,G7864,G7748);
  nand GNAME8072(G8072,G7865,G7972);
  nand GNAME8073(G8073,G7950,G7951,G7952);
  nand GNAME8074(G8074,G7866,G7973);
  nand GNAME8075(G8075,G7946,G7947,G7948);
  nand GNAME8076(G8076,G7867,G7974);
  nand GNAME8077(G8077,G7942,G7943,G7944);
  nand GNAME8078(G8078,G7868,G7975);
  nand GNAME8079(G8079,G7938,G7939,G7940);
  nand GNAME8080(G8080,G7869,G7976);
  nand GNAME8081(G8081,G7912,G7886,G7887);
  nand GNAME8082(G8082,G7870,G7977);
  nand GNAME8083(G8083,G7934,G7935,G7936);
  nand GNAME8084(G8084,G7871,G7978);
  nand GNAME8085(G8085,G7930,G7931,G7932);
  nand GNAME8086(G8086,G7872,G7979);
  nand GNAME8087(G8087,G7926,G7927,G7928);
  nand GNAME8088(G8088,G7725,G7980);
  nand GNAME8089(G8089,G7922,G7923,G7924);
  nand GNAME8090(G8090,G7804,G7751);
  nand GNAME8091(G8091,G7724,G7755);
  nand GNAME8092(G8092,G7723,G7758);
  nand GNAME8093(G8093,G7873,G1278);
  nand GNAME8094(G8094,G7782,G7969);
  not GNAME8095(G8095,G7878);
  not GNAME8096(G8096,G7884);
  not GNAME8097(G8097,G7767);
  not GNAME8098(G8098,G7879);
  not GNAME8099(G8099,G7801);
  not GNAME8100(G8100,G7885);
  nor GNAME8101(G8101,G8105,G8132);
  nor GNAME8102(G8102,G8153,G8107);
  nor GNAME8103(G8103,G8102,G2545);
  and GNAME8104(G8104,G8107,G8153);
  nor GNAME8105(G8105,G8104,G8103,G8151,G8149);
  not GNAME8106(G8106,G2608);
  and GNAME8107(G8107,G8110,G8111);
  not GNAME8108(G8108,G8133);
  nand GNAME8109(G8109,G8106,G8143);
  nand GNAME8110(G8110,G2312,G8108,G8109);
  or GNAME8111(G8111,G8143,G8106);
  or GNAME8112(G8112,G1755,G8113);
  nor GNAME8113(G8113,G557,G556);
  and GNAME8114(G8114,G8130,G8131);
  not GNAME8115(G8115,G21565);
  not GNAME8116(G8116,G1757);
  not GNAME8117(G8117,G21563);
  not GNAME8118(G8118,G1755);
  not GNAME8119(G8119,G1759);
  nand GNAME8120(G8120,G8115,G1758);
  nand GNAME8121(G8121,G21566,G8119,G8120);
  or GNAME8122(G8122,G1758,G8115);
  nand GNAME8123(G8123,G8116,G21564);
  nand GNAME8124(G8124,G8123,G8121,G8122);
  or GNAME8125(G8125,G21564,G8116);
  nand GNAME8126(G8126,G8117,G1756);
  nand GNAME8127(G8127,G8126,G8124,G8125);
  or GNAME8128(G8128,G1756,G8117);
  nand GNAME8129(G8129,G8118,G21562);
  nand GNAME8130(G8130,G8129,G8127,G8128);
  or GNAME8131(G8131,G21562,G8118);
  nand GNAME8132(G8132,G8164,G8167);
  nand GNAME8133(G8133,G8165,G8135);
  not GNAME8134(G8134,G21561);
  or GNAME8135(G8135,G21566,G8134);
  not GNAME8136(G8136,G21560);
  not GNAME8137(G8137,G21564);
  not GNAME8138(G8138,G21559);
  not GNAME8139(G8139,G21563);
  not GNAME8140(G8140,G21558);
  not GNAME8141(G8141,G21562);
  not GNAME8142(G8142,G21557);
  nand GNAME8143(G8143,G8180,G8181);
  and GNAME8144(G8144,G8166,G8167);
  and GNAME8145(G8145,G8170,G8171);
  and GNAME8146(G8146,G8174,G8175);
  and GNAME8147(G8147,G8178,G8179);
  and GNAME8148(G8148,G8162,G8171);
  and GNAME8149(G8149,G8168,G8169);
  and GNAME8150(G8150,G8160,G8175);
  and GNAME8151(G8151,G8172,G8173);
  and GNAME8152(G8152,G8157,G8158);
  and GNAME8153(G8153,G8176,G8177);
  not GNAME8154(G8154,G21565);
  not GNAME8155(G8155,G8135);
  nand GNAME8156(G8156,G8135,G8136);
  nand GNAME8157(G8157,G8154,G8156);
  nand GNAME8158(G8158,G8155,G21560);
  and GNAME8159(G8159,G8138,G21564);
  or GNAME8160(G8160,G8152,G8159);
  and GNAME8161(G8161,G8140,G21563);
  or GNAME8162(G8162,G8150,G8161);
  and GNAME8163(G8163,G8142,G21562);
  or GNAME8164(G8164,G8148,G8163);
  nand GNAME8165(G8165,G8134,G21566);
  nand GNAME8166(G8166,G8142,G21562);
  nand GNAME8167(G8167,G8141,G21557);
  nand GNAME8168(G8168,G8144,G8148);
  or GNAME8169(G8169,G8148,G8144);
  nand GNAME8170(G8170,G8140,G21563);
  nand GNAME8171(G8171,G8139,G21558);
  nand GNAME8172(G8172,G8145,G8150);
  or GNAME8173(G8173,G8150,G8145);
  nand GNAME8174(G8174,G8138,G21564);
  nand GNAME8175(G8175,G8137,G21559);
  nand GNAME8176(G8176,G8146,G8152);
  or GNAME8177(G8177,G8152,G8146);
  nand GNAME8178(G8178,G8136,G21565);
  nand GNAME8179(G8179,G8154,G21560);
  nand GNAME8180(G8180,G8155,G8147);
  or GNAME8181(G8181,G8155,G8147);
  nand GNAME8182(G8182,G8421,G8214);
  and GNAME8183(G8183,G8227,G8214);
  nand GNAME8184(G8184,G8247,G8214);
  nand GNAME8185(G8185,G8246,G8214);
  nand GNAME8186(G8186,G8245,G8214);
  nand GNAME8187(G8187,G8244,G8214);
  nand GNAME8188(G8188,G8243,G8214);
  nand GNAME8189(G8189,G8242,G8214);
  nand GNAME8190(G8190,G8241,G8214);
  nand GNAME8191(G8191,G8240,G8214);
  nand GNAME8192(G8192,G8239,G8214);
  nand GNAME8193(G8193,G8238,G8214);
  nand GNAME8194(G8194,G8237,G8214);
  nand GNAME8195(G8195,G8236,G8214);
  nand GNAME8196(G8196,G8235,G8214);
  nand GNAME8197(G8197,G8234,G8214);
  nand GNAME8198(G8198,G8233,G8214);
  and GNAME8199(G8199,G8232,G8214);
  nand GNAME8200(G8200,G8231,G8214);
  nand GNAME8201(G8201,G8230,G8214);
  nand GNAME8202(G8202,G8229,G8214);
  and GNAME8203(G8203,G8228,G8214);
  nand GNAME8204(G8204,G8224,G8214);
  and GNAME8205(G8205,G8437,G8438);
  and GNAME8206(G8206,G8433,G8435);
  and GNAME8207(G8207,G8429,G8430);
  and GNAME8208(G8208,G8426,G8427);
  and GNAME8209(G8209,G8422,G8424);
  and GNAME8210(G8210,G8420,G8182);
  and GNAME8211(G8211,G8353,G8355);
  and GNAME8212(G8212,G8347,G8348);
  and GNAME8213(G8213,G8343,G8345);
  not GNAME8214(G8214,G1661);
  not GNAME8215(G8215,G724);
  not GNAME8216(G8216,G723);
  not GNAME8217(G8217,G722);
  not GNAME8218(G8218,G721);
  not GNAME8219(G8219,G720);
  not GNAME8220(G8220,G719);
  not GNAME8221(G8221,G718);
  not GNAME8222(G8222,G717);
  not GNAME8223(G8223,G716);
  not GNAME8224(G8224,G715);
  and GNAME8225(G8225,G8341,G8317);
  or GNAME8226(G8226,G8314,G8225);
  not GNAME8227(G8227,G694);
  not GNAME8228(G8228,G714);
  not GNAME8229(G8229,G713);
  not GNAME8230(G8230,G712);
  not GNAME8231(G8231,G711);
  not GNAME8232(G8232,G710);
  not GNAME8233(G8233,G709);
  not GNAME8234(G8234,G708);
  not GNAME8235(G8235,G707);
  not GNAME8236(G8236,G706);
  not GNAME8237(G8237,G705);
  not GNAME8238(G8238,G704);
  not GNAME8239(G8239,G703);
  not GNAME8240(G8240,G702);
  not GNAME8241(G8241,G701);
  not GNAME8242(G8242,G700);
  not GNAME8243(G8243,G699);
  not GNAME8244(G8244,G698);
  not GNAME8245(G8245,G697);
  not GNAME8246(G8246,G696);
  not GNAME8247(G8247,G695);
  nor GNAME8248(G8248,G8183,G8249);
  and GNAME8249(G8249,G8416,G8415);
  and GNAME8250(G8250,G8351,G8323);
  or GNAME8251(G8251,G8320,G8250);
  and GNAME8252(G8252,G8372,G8371);
  nor GNAME8253(G8253,G8199,G8252);
  and GNAME8254(G8254,G8431,G8338);
  or GNAME8255(G8255,G8203,G8254);
  and GNAME8256(G8256,G8474,G8475);
  and GNAME8257(G8257,G8479,G8480);
  nand GNAME8258(G8258,G8528,G8529);
  nand GNAME8259(G8259,G8484,G8485);
  nand GNAME8260(G8260,G8486,G8487);
  nand GNAME8261(G8261,G8488,G8489);
  nand GNAME8262(G8262,G8490,G8491);
  nand GNAME8263(G8263,G8492,G8493);
  nand GNAME8264(G8264,G8494,G8495);
  nand GNAME8265(G8265,G8496,G8497);
  nand GNAME8266(G8266,G8498,G8499);
  nand GNAME8267(G8267,G8500,G8501);
  nand GNAME8268(G8268,G8502,G8503);
  nand GNAME8269(G8269,G8504,G8505);
  nand GNAME8270(G8270,G8506,G8507);
  nand GNAME8271(G8271,G8508,G8509);
  nand GNAME8272(G8272,G8510,G8511);
  nand GNAME8273(G8273,G8512,G8513);
  nand GNAME8274(G8274,G8514,G8515);
  nand GNAME8275(G8275,G8516,G8517);
  nand GNAME8276(G8276,G8518,G8519);
  nand GNAME8277(G8277,G8520,G8521);
  nand GNAME8278(G8278,G8522,G8523);
  nand GNAME8279(G8279,G8524,G8525);
  nand GNAME8280(G8280,G8526,G8527);
  not GNAME8281(G8281,G685);
  not GNAME8282(G8282,G686);
  not GNAME8283(G8283,G687);
  not GNAME8284(G8284,G689);
  not GNAME8285(G8285,G690);
  not GNAME8286(G8286,G691);
  nand GNAME8287(G8287,G8334,G8313);
  nand GNAME8288(G8288,G8339,G8311);
  nand GNAME8289(G8289,G8328,G8319);
  nand GNAME8290(G8290,G8413,G8412);
  nand GNAME8291(G8291,G8410,G8409);
  nand GNAME8292(G8292,G8407,G8406);
  nand GNAME8293(G8293,G8404,G8403);
  nand GNAME8294(G8294,G8401,G8400);
  nand GNAME8295(G8295,G8398,G8397);
  nand GNAME8296(G8296,G8395,G8394);
  nand GNAME8297(G8297,G8392,G8391);
  nand GNAME8298(G8298,G8389,G8388);
  nand GNAME8299(G8299,G8386,G8385);
  nand GNAME8300(G8300,G8349,G8310);
  nand GNAME8301(G8301,G8383,G8382);
  nand GNAME8302(G8302,G8380,G8379);
  nand GNAME8303(G8303,G8377,G8376);
  nand GNAME8304(G8304,G8374,G8357);
  or GNAME8305(G8305,G8253,G8358);
  nand GNAME8306(G8306,G8369,G8368);
  nand GNAME8307(G8307,G8366,G8359);
  nand GNAME8308(G8308,G8324,G8310);
  or GNAME8309(G8309,G8214,G8223);
  or GNAME8310(G8310,G8256,G8215);
  or GNAME8311(G8311,G8257,G8219);
  nand GNAME8312(G8312,G8222,G8462,G8463);
  nand GNAME8313(G8313,G8483,G717);
  and GNAME8314(G8314,G8221,G8464,G8465);
  nand GNAME8315(G8315,G8482,G718);
  nand GNAME8316(G8316,G8220,G8466,G8467);
  nand GNAME8317(G8317,G8481,G719);
  nand GNAME8318(G8318,G8218,G8468,G8469);
  nand GNAME8319(G8319,G8478,G721);
  and GNAME8320(G8320,G8217,G8470,G8471);
  nand GNAME8321(G8321,G8477,G722);
  nand GNAME8322(G8322,G8216,G8472,G8473);
  nand GNAME8323(G8323,G8476,G723);
  nand GNAME8324(G8324,G8215,G8256);
  nand GNAME8325(G8325,G8351,G8323);
  nand GNAME8326(G8326,G8531,G8325);
  nand GNAME8327(G8327,G8326,G8321);
  nand GNAME8328(G8328,G8318,G8327);
  not GNAME8329(G8329,G8289);
  nand GNAME8330(G8330,G8219,G8257);
  nand GNAME8331(G8331,G8341,G8317);
  nand GNAME8332(G8332,G8530,G8331);
  nand GNAME8333(G8333,G8332,G8315);
  nand GNAME8334(G8334,G8312,G8333);
  not GNAME8335(G8335,G8287);
  nand GNAME8336(G8336,G8223,G8214);
  not GNAME8337(G8337,G8362);
  nand GNAME8338(G8338,G1661,G715);
  nand GNAME8339(G8339,G8289,G8330);
  not GNAME8340(G8340,G8288);
  nand GNAME8341(G8341,G8316,G8288);
  nand GNAME8342(G8342,G8315,G8226);
  nand GNAME8343(G8343,G8342,G8312,G8313);
  nand GNAME8344(G8344,G8312,G8313);
  nand GNAME8345(G8345,G8344,G8315,G8226);
  or GNAME8346(G8346,G8314,G8533);
  nand GNAME8347(G8347,G8346,G8225);
  or GNAME8348(G8348,G8533,G8226);
  nand GNAME8349(G8349,G8324,G1661);
  not GNAME8350(G8350,G8300);
  nand GNAME8351(G8351,G8322,G8300);
  nand GNAME8352(G8352,G8321,G8251);
  nand GNAME8353(G8353,G8352,G8318,G8319);
  nand GNAME8354(G8354,G8318,G8319);
  nand GNAME8355(G8355,G8354,G8321,G8251);
  and GNAME8356(G8356,G1661,G694);
  nand GNAME8357(G8357,G1661,G709);
  and GNAME8358(G8358,G1661,G710);
  nand GNAME8359(G8359,G1661,G713);
  nand GNAME8360(G8360,G1661,G714);
  nand GNAME8361(G8361,G8287,G8336);
  nand GNAME8362(G8362,G8361,G8309);
  nand GNAME8363(G8363,G8431,G8338);
  nand GNAME8364(G8364,G8532,G8363);
  nand GNAME8365(G8365,G8364,G8360);
  nand GNAME8366(G8366,G8202,G8365);
  not GNAME8367(G8367,G8307);
  nand GNAME8368(G8368,G1661,G712);
  nand GNAME8369(G8369,G8307,G8201);
  not GNAME8370(G8370,G8306);
  nand GNAME8371(G8371,G1661,G711);
  nand GNAME8372(G8372,G8306,G8200);
  not GNAME8373(G8373,G8305);
  nand GNAME8374(G8374,G8198,G8305);
  not GNAME8375(G8375,G8304);
  nand GNAME8376(G8376,G1661,G708);
  nand GNAME8377(G8377,G8304,G8197);
  not GNAME8378(G8378,G8303);
  nand GNAME8379(G8379,G1661,G707);
  nand GNAME8380(G8380,G8303,G8196);
  not GNAME8381(G8381,G8302);
  nand GNAME8382(G8382,G1661,G706);
  nand GNAME8383(G8383,G8302,G8195);
  not GNAME8384(G8384,G8301);
  nand GNAME8385(G8385,G1661,G705);
  nand GNAME8386(G8386,G8301,G8194);
  not GNAME8387(G8387,G8299);
  nand GNAME8388(G8388,G1661,G704);
  nand GNAME8389(G8389,G8299,G8193);
  not GNAME8390(G8390,G8298);
  nand GNAME8391(G8391,G1661,G703);
  nand GNAME8392(G8392,G8298,G8192);
  not GNAME8393(G8393,G8297);
  nand GNAME8394(G8394,G1661,G702);
  nand GNAME8395(G8395,G8297,G8191);
  not GNAME8396(G8396,G8296);
  nand GNAME8397(G8397,G1661,G701);
  nand GNAME8398(G8398,G8296,G8190);
  not GNAME8399(G8399,G8295);
  nand GNAME8400(G8400,G1661,G700);
  nand GNAME8401(G8401,G8295,G8189);
  not GNAME8402(G8402,G8294);
  nand GNAME8403(G8403,G1661,G699);
  nand GNAME8404(G8404,G8294,G8188);
  not GNAME8405(G8405,G8293);
  nand GNAME8406(G8406,G1661,G698);
  nand GNAME8407(G8407,G8293,G8187);
  not GNAME8408(G8408,G8292);
  nand GNAME8409(G8409,G1661,G697);
  nand GNAME8410(G8410,G8292,G8186);
  not GNAME8411(G8411,G8291);
  nand GNAME8412(G8412,G1661,G696);
  nand GNAME8413(G8413,G8291,G8185);
  not GNAME8414(G8414,G8290);
  nand GNAME8415(G8415,G1661,G695);
  nand GNAME8416(G8416,G8290,G8184);
  or GNAME8417(G8417,G8356,G8248);
  nand GNAME8418(G8418,G8417,G693);
  or GNAME8419(G8419,G8248,G693,G8356);
  nand GNAME8420(G8420,G1661,G8418,G8419);
  nand GNAME8421(G8421,G8418,G8419);
  or GNAME8422(G8422,G8356,G8534);
  or GNAME8423(G8423,G8356,G8183);
  nand GNAME8424(G8424,G8423,G8249);
  or GNAME8425(G8425,G8320,G8535);
  nand GNAME8426(G8426,G8425,G8250);
  or GNAME8427(G8427,G8535,G8251);
  or GNAME8428(G8428,G8358,G8199);
  nand GNAME8429(G8429,G8428,G8252);
  or GNAME8430(G8430,G8358,G8536);
  nand GNAME8431(G8431,G8362,G8204);
  nand GNAME8432(G8432,G8360,G8255);
  nand GNAME8433(G8433,G8432,G8202,G8359);
  nand GNAME8434(G8434,G8202,G8359);
  nand GNAME8435(G8435,G8434,G8360,G8255);
  or GNAME8436(G8436,G8203,G8537);
  nand GNAME8437(G8437,G8436,G8254);
  or GNAME8438(G8438,G8537,G8255);
  not GNAME8439(G8439,G8308);
  nand GNAME8440(G8440,G8204,G8338);
  nand GNAME8441(G8441,G8309,G8336);
  nand GNAME8442(G8442,G8316,G8317);
  nand GNAME8443(G8443,G8311,G8330);
  nand GNAME8444(G8444,G8184,G8415);
  nand GNAME8445(G8445,G8185,G8412);
  nand GNAME8446(G8446,G8186,G8409);
  nand GNAME8447(G8447,G8187,G8406);
  nand GNAME8448(G8448,G8188,G8403);
  nand GNAME8449(G8449,G8189,G8400);
  nand GNAME8450(G8450,G8190,G8397);
  nand GNAME8451(G8451,G8191,G8394);
  nand GNAME8452(G8452,G8192,G8391);
  nand GNAME8453(G8453,G8193,G8388);
  nand GNAME8454(G8454,G8322,G8323);
  nand GNAME8455(G8455,G8194,G8385);
  nand GNAME8456(G8456,G8195,G8382);
  nand GNAME8457(G8457,G8196,G8379);
  nand GNAME8458(G8458,G8197,G8376);
  nand GNAME8459(G8459,G8198,G8357);
  nand GNAME8460(G8460,G8200,G8371);
  nand GNAME8461(G8461,G8201,G8368);
  nand GNAME8462(G8462,G8281,G1661);
  nand GNAME8463(G8463,G8214,G685);
  nand GNAME8464(G8464,G8282,G1661);
  nand GNAME8465(G8465,G8214,G686);
  nand GNAME8466(G8466,G8283,G1661);
  nand GNAME8467(G8467,G8214,G687);
  nand GNAME8468(G8468,G8284,G1661);
  nand GNAME8469(G8469,G8214,G689);
  nand GNAME8470(G8470,G8285,G1661);
  nand GNAME8471(G8471,G8214,G690);
  nand GNAME8472(G8472,G8286,G1661);
  nand GNAME8473(G8473,G8214,G691);
  or GNAME8474(G8474,G692,G8214);
  nand GNAME8475(G8475,G8214,G692);
  nand GNAME8476(G8476,G8472,G8473);
  nand GNAME8477(G8477,G8470,G8471);
  nand GNAME8478(G8478,G8468,G8469);
  or GNAME8479(G8479,G688,G8214);
  nand GNAME8480(G8480,G8214,G688);
  nand GNAME8481(G8481,G8466,G8467);
  nand GNAME8482(G8482,G8464,G8465);
  nand GNAME8483(G8483,G8462,G8463);
  nand GNAME8484(G8484,G8362,G8440);
  nand GNAME8485(G8485,G8337,G8204,G8338);
  nand GNAME8486(G8486,G8287,G8441);
  nand GNAME8487(G8487,G8335,G8309,G8336);
  nand GNAME8488(G8488,G8288,G8442);
  nand GNAME8489(G8489,G8340,G8316,G8317);
  nand GNAME8490(G8490,G8289,G8443);
  nand GNAME8491(G8491,G8329,G8311,G8330);
  nand GNAME8492(G8492,G8290,G8444);
  nand GNAME8493(G8493,G8414,G8184,G8415);
  nand GNAME8494(G8494,G8291,G8445);
  nand GNAME8495(G8495,G8411,G8185,G8412);
  nand GNAME8496(G8496,G8292,G8446);
  nand GNAME8497(G8497,G8408,G8186,G8409);
  nand GNAME8498(G8498,G8293,G8447);
  nand GNAME8499(G8499,G8405,G8187,G8406);
  nand GNAME8500(G8500,G8294,G8448);
  nand GNAME8501(G8501,G8402,G8188,G8403);
  nand GNAME8502(G8502,G8295,G8449);
  nand GNAME8503(G8503,G8399,G8189,G8400);
  nand GNAME8504(G8504,G8296,G8450);
  nand GNAME8505(G8505,G8396,G8190,G8397);
  nand GNAME8506(G8506,G8297,G8451);
  nand GNAME8507(G8507,G8393,G8191,G8394);
  nand GNAME8508(G8508,G8298,G8452);
  nand GNAME8509(G8509,G8390,G8192,G8391);
  nand GNAME8510(G8510,G8299,G8453);
  nand GNAME8511(G8511,G8387,G8193,G8388);
  nand GNAME8512(G8512,G8300,G8454);
  nand GNAME8513(G8513,G8350,G8322,G8323);
  nand GNAME8514(G8514,G8301,G8455);
  nand GNAME8515(G8515,G8384,G8194,G8385);
  nand GNAME8516(G8516,G8302,G8456);
  nand GNAME8517(G8517,G8381,G8195,G8382);
  nand GNAME8518(G8518,G8303,G8457);
  nand GNAME8519(G8519,G8378,G8196,G8379);
  nand GNAME8520(G8520,G8304,G8458);
  nand GNAME8521(G8521,G8375,G8197,G8376);
  nand GNAME8522(G8522,G8305,G8459);
  nand GNAME8523(G8523,G8373,G8198,G8357);
  nand GNAME8524(G8524,G8306,G8460);
  nand GNAME8525(G8525,G8370,G8200,G8371);
  nand GNAME8526(G8526,G8307,G8461);
  nand GNAME8527(G8527,G8367,G8201,G8368);
  nand GNAME8528(G8528,G8308,G1661);
  nand GNAME8529(G8529,G8214,G8439);
  not GNAME8530(G8530,G8314);
  not GNAME8531(G8531,G8320);
  not GNAME8532(G8532,G8203);
  not GNAME8533(G8533,G8315);
  not GNAME8534(G8534,G8248);
  not GNAME8535(G8535,G8321);
  not GNAME8536(G8536,G8253);
  not GNAME8537(G8537,G8360);
  and GNAME8538(G8538,G8633,G8634);
  nand GNAME8539(G8539,G8635,G8639,G8640);
  not GNAME8540(G8540,G7811);
  nand GNAME8541(G8541,G575,G7811);
  not GNAME8542(G8542,G7810);
  not GNAME8543(G8543,G7773);
  not GNAME8544(G8544,G573);
  not GNAME8545(G8545,G7774);
  not GNAME8546(G8546,G572);
  not GNAME8547(G8547,G7831);
  not GNAME8548(G8548,G571);
  not GNAME8549(G8549,G7830);
  not GNAME8550(G8550,G570);
  not GNAME8551(G8551,G7775);
  not GNAME8552(G8552,G569);
  not GNAME8553(G8553,G7827);
  not GNAME8554(G8554,G7828);
  nor GNAME8555(G8555,G8554,G8603,G8553);
  not GNAME8556(G8556,G7826);
  and GNAME8557(G8557,G8555,G7826);
  not GNAME8558(G8558,G7825);
  and GNAME8559(G8559,G8557,G7825);
  not GNAME8560(G8560,G7823);
  and GNAME8561(G8561,G8559,G7823);
  not GNAME8562(G8562,G7822);
  and GNAME8563(G8563,G8561,G7822);
  not GNAME8564(G8564,G7821);
  and GNAME8565(G8565,G8563,G7821);
  not GNAME8566(G8566,G7820);
  and GNAME8567(G8567,G8565,G7820);
  not GNAME8568(G8568,G7819);
  and GNAME8569(G8569,G8567,G7819);
  not GNAME8570(G8570,G7818);
  and GNAME8571(G8571,G8569,G7818);
  not GNAME8572(G8572,G7817);
  and GNAME8573(G8573,G8571,G7817);
  not GNAME8574(G8574,G7816);
  not GNAME8575(G8575,G7815);
  nand GNAME8576(G8576,G7815,G8573,G7816);
  and GNAME8577(G8577,G8628,G8629);
  nor GNAME8578(G8578,G8630,G8577);
  nand GNAME8579(G8579,G8641,G8642);
  nand GNAME8580(G8580,G8643,G8644);
  nand GNAME8581(G8581,G8645,G8646);
  nand GNAME8582(G8582,G8647,G8648);
  nand GNAME8583(G8583,G8649,G8650);
  nand GNAME8584(G8584,G8651,G8652);
  nand GNAME8585(G8585,G8653,G8654);
  nand GNAME8586(G8586,G8655,G8656);
  nand GNAME8587(G8587,G8657,G8658);
  nand GNAME8588(G8588,G8659,G8660);
  nand GNAME8589(G8589,G8661,G8662);
  nand GNAME8590(G8590,G8663,G8664);
  nand GNAME8591(G8591,G8665,G8666);
  nand GNAME8592(G8592,G8667,G8668);
  nand GNAME8593(G8593,G8669,G8670);
  nand GNAME8594(G8594,G8676,G8677);
  nand GNAME8595(G8595,G8681,G8682);
  nand GNAME8596(G8596,G8686,G8687);
  nand GNAME8597(G8597,G8691,G8692);
  nand GNAME8598(G8598,G8696,G8697);
  nand GNAME8599(G8599,G8611,G574);
  nand GNAME8600(G8600,G7814,G8699);
  and GNAME8601(G8601,G8573,G7816);
  nor GNAME8602(G8602,G8603,G8554);
  nor GNAME8603(G8603,G8698,G8578);
  and GNAME8604(G8604,G8671,G8672);
  nand GNAME8605(G8605,G8625,G8626);
  nand GNAME8606(G8606,G8622,G8623);
  nand GNAME8607(G8607,G8619,G8620);
  nand GNAME8608(G8608,G8616,G8617);
  nand GNAME8609(G8609,G8614,G8599);
  not GNAME8610(G8610,G8603);
  not GNAME8611(G8611,G8541);
  nand GNAME8612(G8612,G7829,G568);
  or GNAME8613(G8613,G8611,G574);
  nand GNAME8614(G8614,G8613,G7810);
  nand GNAME8615(G8615,G8544,G8543);
  nand GNAME8616(G8616,G8609,G8615);
  or GNAME8617(G8617,G8543,G8544);
  nand GNAME8618(G8618,G8546,G8545);
  nand GNAME8619(G8619,G8608,G8618);
  or GNAME8620(G8620,G8545,G8546);
  nand GNAME8621(G8621,G8548,G8547);
  nand GNAME8622(G8622,G8607,G8621);
  or GNAME8623(G8623,G8547,G8548);
  nand GNAME8624(G8624,G8550,G8549);
  nand GNAME8625(G8625,G8606,G8624);
  or GNAME8626(G8626,G8549,G8550);
  nand GNAME8627(G8627,G8552,G8551);
  nand GNAME8628(G8628,G8605,G8627);
  or GNAME8629(G8629,G8551,G8552);
  nor GNAME8630(G8630,G7829,G568);
  or GNAME8631(G8631,G568,G7829);
  nand GNAME8632(G8632,G8612,G8631);
  nand GNAME8633(G8633,G8632,G8577);
  nand GNAME8634(G8634,G8612,G8578);
  or GNAME8635(G8635,G574,G8638);
  or GNAME8636(G8636,G8611,G8542);
  or GNAME8637(G8637,G7810,G8541);
  and GNAME8638(G8638,G8636,G8637);
  nand GNAME8639(G8639,G8542,G8541,G574);
  or GNAME8640(G8640,G8542,G8599);
  or GNAME8641(G8641,G575,G8540);
  nand GNAME8642(G8642,G8540,G575);
  nand GNAME8643(G8643,G8600,G7777);
  or GNAME8644(G8644,G7777,G8600);
  or GNAME8645(G8645,G7814,G8576);
  nand GNAME8646(G8646,G8576,G7814);
  or GNAME8647(G8647,G8601,G8575);
  nand GNAME8648(G8648,G8575,G8601);
  or GNAME8649(G8649,G8573,G8574);
  nand GNAME8650(G8650,G8574,G8573);
  or GNAME8651(G8651,G8571,G8572);
  nand GNAME8652(G8652,G8572,G8571);
  or GNAME8653(G8653,G8569,G8570);
  nand GNAME8654(G8654,G8570,G8569);
  or GNAME8655(G8655,G8567,G8568);
  nand GNAME8656(G8656,G8568,G8567);
  or GNAME8657(G8657,G8565,G8566);
  nand GNAME8658(G8658,G8566,G8565);
  or GNAME8659(G8659,G8563,G8564);
  nand GNAME8660(G8660,G8564,G8563);
  or GNAME8661(G8661,G8561,G8562);
  nand GNAME8662(G8662,G8562,G8561);
  or GNAME8663(G8663,G8559,G8560);
  nand GNAME8664(G8664,G8560,G8559);
  or GNAME8665(G8665,G8557,G8558);
  nand GNAME8666(G8666,G8558,G8557);
  or GNAME8667(G8667,G8555,G8556);
  nand GNAME8668(G8668,G8556,G8555);
  or GNAME8669(G8669,G8602,G8553);
  nand GNAME8670(G8670,G8553,G8602);
  or GNAME8671(G8671,G8603,G8554);
  or GNAME8672(G8672,G7828,G8610);
  or GNAME8673(G8673,G7775,G8552);
  or GNAME8674(G8674,G569,G8551);
  and GNAME8675(G8675,G8673,G8674);
  nand GNAME8676(G8676,G8605,G8673,G8674);
  or GNAME8677(G8677,G8675,G8605);
  or GNAME8678(G8678,G7830,G8550);
  or GNAME8679(G8679,G570,G8549);
  and GNAME8680(G8680,G8678,G8679);
  nand GNAME8681(G8681,G8606,G8678,G8679);
  or GNAME8682(G8682,G8680,G8606);
  or GNAME8683(G8683,G7831,G8548);
  or GNAME8684(G8684,G571,G8547);
  and GNAME8685(G8685,G8683,G8684);
  nand GNAME8686(G8686,G8607,G8683,G8684);
  or GNAME8687(G8687,G8685,G8607);
  or GNAME8688(G8688,G7774,G8546);
  or GNAME8689(G8689,G572,G8545);
  and GNAME8690(G8690,G8688,G8689);
  nand GNAME8691(G8691,G8608,G8688,G8689);
  or GNAME8692(G8692,G8690,G8608);
  or GNAME8693(G8693,G7773,G8544);
  or GNAME8694(G8694,G573,G8543);
  and GNAME8695(G8695,G8693,G8694);
  nand GNAME8696(G8696,G8609,G8693,G8694);
  or GNAME8697(G8697,G8695,G8609);
  not GNAME8698(G8698,G8612);
  not GNAME8699(G8699,G8576);
  not GNAME8700(G8700,G1753);
  not GNAME8701(G8701,G1754);
  not GNAME8702(G8702,G559);
  not GNAME8703(G8703,G1752);
  nor GNAME8704(G8704,G8749,G8831);
  and GNAME8705(G8705,G8825,G8829);
  nor GNAME8706(G8706,G8751,G8828);
  and GNAME8707(G8707,G8752,G8826);
  nand GNAME8708(G8708,G8834,G8856,G8857);
  and GNAME8709(G8709,G8710,G8832);
  nand GNAME8710(G8710,G2511,G748);
  not GNAME8711(G8711,G747);
  and GNAME8712(G8712,G8797,G747);
  not GNAME8713(G8713,G2511);
  not GNAME8714(G8714,G745);
  and GNAME8715(G8715,G8781,G745);
  not GNAME8716(G8716,G743);
  not GNAME8717(G8717,G744);
  not GNAME8718(G8718,G741);
  and GNAME8719(G8719,G744,G8715,G743);
  not GNAME8720(G8720,G742);
  and GNAME8721(G8721,G742,G741,G8719);
  not GNAME8722(G8722,G740);
  and GNAME8723(G8723,G8721,G740);
  and GNAME8724(G8724,G739,G8723);
  not GNAME8725(G8725,G737);
  not GNAME8726(G8726,G738);
  not GNAME8727(G8727,G735);
  and GNAME8728(G8728,G738,G8724,G737);
  not GNAME8729(G8729,G736);
  not GNAME8730(G8730,G733);
  and GNAME8731(G8731,G736,G735,G8728);
  not GNAME8732(G8732,G734);
  and GNAME8733(G8733,G734,G733,G8731);
  not GNAME8734(G8734,G732);
  not GNAME8735(G8735,G731);
  not GNAME8736(G8736,G755);
  not GNAME8737(G8737,G730);
  not GNAME8738(G8738,G754);
  not GNAME8739(G8739,G729);
  not GNAME8740(G8740,G753);
  not GNAME8741(G8741,G728);
  not GNAME8742(G8742,G752);
  not GNAME8743(G8743,G727);
  not GNAME8744(G8744,G751);
  not GNAME8745(G8745,G726);
  not GNAME8746(G8746,G750);
  not GNAME8747(G8747,G1768);
  not GNAME8748(G8748,G749);
  and GNAME8749(G8749,G1767,G8784,G1766);
  and GNAME8750(G8750,G8749,G1765);
  and GNAME8751(G8751,G1764,G8750,G1763);
  nand GNAME8752(G8752,G8751,G1762);
  not GNAME8753(G8753,G1761);
  nand GNAME8754(G8754,G8835,G8836);
  nand GNAME8755(G8755,G8837,G8838);
  nand GNAME8756(G8756,G8839,G8840);
  nand GNAME8757(G8757,G8841,G8842);
  nand GNAME8758(G8758,G8843,G8844);
  nand GNAME8759(G8759,G8845,G8846);
  nand GNAME8760(G8760,G8851,G8852);
  nand GNAME8761(G8761,G8858,G8859);
  nand GNAME8762(G8762,G8882,G8883);
  nand GNAME8763(G8763,G7312,G7311);
  nand GNAME8764(G8764,G7310,G7309);
  nand GNAME8765(G8765,G7308,G7307);
  nand GNAME8766(G8766,G7306,G7305);
  nand GNAME8767(G8767,G7304,G7303);
  nand GNAME8768(G8768,G7302,G7301);
  nand GNAME8769(G8769,G7300,G7299);
  nand GNAME8770(G8770,G8849,G8850);
  nand GNAME8771(G8771,G8865,G8866);
  nand GNAME8772(G8772,G8870,G8871);
  nand GNAME8773(G8773,G8875,G8876);
  nand GNAME8774(G8774,G8880,G8881);
  nand GNAME8775(G8775,G8887,G8888);
  nand GNAME8776(G8776,G8892,G8893);
  nand GNAME8777(G8777,G7316,G7315);
  and GNAME8778(G8778,G7314,G7313);
  and GNAME8779(G8779,G8719,G742);
  and GNAME8780(G8780,G8715,G744);
  or GNAME8781(G8781,G8799,G8783);
  and GNAME8782(G8782,G8847,G8848);
  and GNAME8783(G8783,G8712,G2511);
  nand GNAME8784(G8784,G8823,G8824);
  and GNAME8785(G8785,G8860,G8861);
  nand GNAME8786(G8786,G8820,G8821);
  nand GNAME8787(G8787,G8817,G8818);
  nand GNAME8788(G8788,G8814,G8815);
  nand GNAME8789(G8789,G8811,G8812);
  nand GNAME8790(G8790,G8808,G8809);
  nand GNAME8791(G8791,G8805,G8806);
  nand GNAME8792(G8792,G8802,G8803);
  and GNAME8793(G8793,G8731,G734);
  and GNAME8794(G8794,G8728,G736);
  and GNAME8795(G8795,G8724,G738);
  not GNAME8796(G8796,G8712);
  not GNAME8797(G8797,G8710);
  nand GNAME8798(G8798,G8796,G8713);
  and GNAME8799(G8799,G8798,G746);
  not GNAME8800(G8800,G8781);
  or GNAME8801(G8801,G8733,G732);
  nand GNAME8802(G8802,G8801,G756);
  nand GNAME8803(G8803,G8733,G732);
  or GNAME8804(G8804,G755,G731);
  nand GNAME8805(G8805,G8792,G8804);
  nand GNAME8806(G8806,G731,G755);
  or GNAME8807(G8807,G754,G730);
  nand GNAME8808(G8808,G8791,G8807);
  nand GNAME8809(G8809,G730,G754);
  or GNAME8810(G8810,G753,G729);
  nand GNAME8811(G8811,G8790,G8810);
  nand GNAME8812(G8812,G729,G753);
  or GNAME8813(G8813,G752,G728);
  nand GNAME8814(G8814,G8789,G8813);
  nand GNAME8815(G8815,G728,G752);
  or GNAME8816(G8816,G751,G727);
  nand GNAME8817(G8817,G8788,G8816);
  nand GNAME8818(G8818,G727,G751);
  or GNAME8819(G8819,G750,G726);
  nand GNAME8820(G8820,G8787,G8819);
  nand GNAME8821(G8821,G726,G750);
  or GNAME8822(G8822,G749,G1768);
  nand GNAME8823(G8823,G8786,G8822);
  nand GNAME8824(G8824,G1768,G749);
  not GNAME8825(G8825,G8750);
  or GNAME8826(G8826,G8751,G1762);
  and GNAME8827(G8827,G8750,G1764);
  nor GNAME8828(G8828,G8827,G1763);
  or GNAME8829(G8829,G8749,G1765);
  and GNAME8830(G8830,G8784,G1767);
  nor GNAME8831(G8831,G8830,G1766);
  or GNAME8832(G8832,G748,G2511);
  or GNAME8833(G8833,G8752,G8753);
  nand GNAME8834(G8834,G8713,G8855);
  nand GNAME8835(G8835,G7298,G739);
  or GNAME8836(G8836,G739,G7298);
  or GNAME8837(G8837,G8721,G8722);
  nand GNAME8838(G8838,G8722,G8721);
  or GNAME8839(G8839,G8779,G8718);
  nand GNAME8840(G8840,G8718,G8779);
  or GNAME8841(G8841,G8719,G8720);
  nand GNAME8842(G8842,G8720,G8719);
  or GNAME8843(G8843,G8780,G8716);
  nand GNAME8844(G8844,G8716,G8780);
  or GNAME8845(G8845,G8715,G8717);
  nand GNAME8846(G8846,G8717,G8715);
  nand GNAME8847(G8847,G8781,G745);
  nand GNAME8848(G8848,G8714,G8800);
  nand GNAME8849(G8849,G8833,G725);
  or GNAME8850(G8850,G725,G8752,G8753);
  nand GNAME8851(G8851,G8752,G1761);
  or GNAME8852(G8852,G1761,G8752);
  nand GNAME8853(G8853,G8796,G746);
  or GNAME8854(G8854,G746,G8796);
  nand GNAME8855(G8855,G8853,G8854);
  or GNAME8856(G8856,G746,G8712,G8713);
  nand GNAME8857(G8857,G746,G8783);
  nand GNAME8858(G8858,G8825,G1764);
  or GNAME8859(G8859,G1764,G8825);
  nand GNAME8860(G8860,G8784,G1767);
  or GNAME8861(G8861,G1767,G8784);
  nand GNAME8862(G8862,G8747,G749);
  nand GNAME8863(G8863,G8748,G1768);
  and GNAME8864(G8864,G8862,G8863);
  nand GNAME8865(G8865,G8786,G8862,G8863);
  or GNAME8866(G8866,G8864,G8786);
  nand GNAME8867(G8867,G8745,G750);
  nand GNAME8868(G8868,G8746,G726);
  and GNAME8869(G8869,G8867,G8868);
  nand GNAME8870(G8870,G8787,G8867,G8868);
  or GNAME8871(G8871,G8869,G8787);
  nand GNAME8872(G8872,G8743,G751);
  nand GNAME8873(G8873,G8744,G727);
  and GNAME8874(G8874,G8872,G8873);
  nand GNAME8875(G8875,G8788,G8872,G8873);
  or GNAME8876(G8876,G8874,G8788);
  nand GNAME8877(G8877,G8741,G752);
  nand GNAME8878(G8878,G8742,G728);
  and GNAME8879(G8879,G8877,G8878);
  nand GNAME8880(G8880,G8789,G8877,G8878);
  or GNAME8881(G8881,G8879,G8789);
  nand GNAME8882(G8882,G8710,G747);
  nand GNAME8883(G8883,G8711,G8797);
  nand GNAME8884(G8884,G8739,G753);
  nand GNAME8885(G8885,G8740,G729);
  and GNAME8886(G8886,G8884,G8885);
  nand GNAME8887(G8887,G8790,G8884,G8885);
  or GNAME8888(G8888,G8886,G8790);
  nand GNAME8889(G8889,G8737,G754);
  nand GNAME8890(G8890,G8738,G730);
  and GNAME8891(G8891,G8889,G8890);
  nand GNAME8892(G8892,G8791,G8889,G8890);
  or GNAME8893(G8893,G8891,G8791);

endmodule
